//
// Verilog description for cell top, 
// 05/05/15 12:36:35
//
// Precision RTL Plus , 2011a.61//


module top ( CLK, RST, KEY, DATA, READ, STB_DATA, STB_KEY, DATA_OUT, SIGN_REG
              ) ;

    input CLK ;
    input RST ;
    input KEY ;
    input [7:0]DATA ;
    input READ ;
    input STB_DATA ;
    input STB_KEY ;
    output [7:0]DATA_OUT ;
    output [7:0]SIGN_REG ;

    wire [7:2]SIGN_REG_dup_0;
    wire [7:0]STREAM;
    wire WRITE;
    wire [92:0]ENCR_DEV_reg_str_1;
    wire [83:0]ENCR_DEV_reg_str_2;
    wire [110:0]ENCR_DEV_reg_str_3;
    wire [11:0]ENCR_DEV_cnt_init;
    wire [63:0]ENCR_DEV_err_cnt;
    wire [6:0]ENCR_DEV_key_cnt;
    wire [8:0]ENCR_DEV_encry_cnt;
    wire [7:0]ENCR_DEV_data_reg;
    wire [79:0]ENCR_DEV_key_reg;
    wire ENCR_DEV_strob_data_tmp;
    wire [8:0]ENCR_DEV_prev;
    wire [7:0]FIFO_DEV_count;
    wire [0:255]FIFO_DEV_rtlc_msr_n3;
    wire [7:0]FIFO_DEV_rtlc_wadd_n4;
    wire [7:0]FIFO_DEV_rtlc_radd_N1;
    wire nx12521z1, nx12521z6, nx12521z4, nx11524z2, nx10527z2, nx9530z2, 
         nx8533z2, nx7536z2, nx6539z2, nx5542z2, nx12521z11, nx12521z8, 
         nx11524z4, nx10527z4, nx9530z4, nx8533z4, nx7536z4, nx6539z4, nx5542z4, 
         CLK_int, RST_int, KEY_int;
    wire [7:0]DATA_int;
    wire READ_int, STB_DATA_int, STB_KEY_int;
    wire [7:0]DATA_OUT_dup_0;
    wire CONDITION_1_, NOT_CONDITION_0_, ENCR_DEV_t_1_0_, ENCR_DEV_t_1_1_, 
         ENCR_DEV_t_1_2_, ENCR_DEV_t_1_3_, ENCR_DEV_t_1_5_, ENCR_DEV_t_1_6_;
    
    wire [0:7]ENCR_DEV_t_2;
    wire [0:7]ENCR_DEV_t_3;
    wire ENCR_DEV_PWR, nx7516z2, nx3438z3, nx14495z3, nx14495z4, nx14495z2, 
         nx15492z5, nx15492z3;
    wire [79:0]ENCR_DEV_key_reg_12n5ss1;
    wire ENCR_DEV_rtlc12_X_0_n169;
    wire [7:0]ENCR_DEV_stream_15n2ss1;
    wire [92:0]ENCR_DEV_reg_str_1_15n2ss1;
    wire [83:0]ENCR_DEV_reg_str_2_15n2ss1;
    wire [110:0]ENCR_DEV_reg_str_3_15n2ss1;
    wire nx8587z1, nx63528z1, nx46110z1, NOT_ENCR_DEV_t_1_4_16n1s20, 
         NOT_ENCR_DEV_t_1_7_16n1s32, nx18636z1, nx1908z1, nx10507z1, nx9510z1, 
         nx15492z1, nx36622z1, nx13498z1, nx11504z1, nx7516z1, nx14495z1, 
         nx3438z1, nx3438z5, nx10507z5, nx9510z9, nx15492z2, nx36622z3, 
         nx11504z22, nx45632z3, nx25368z1, nx9510z3, nx10507z3, nx35008z1, 
         nx13690z1, nx16127z1, nx37999z1, nx22109z1, nx36005z1, nx21112z1, 
         nx12693z1, nx38996z1, nx37002z1, nx20115z1, nx11696z1, nx39993z1, 
         nx19118z1, nx10699z1, nx40990z1, nx18121z1, nx22484z2, nx41987z1, 
         nx17124z1, nx8705z1, nx7708z1, nx15130z1, nx25475z2, nx12521z5, 
         nx32158z2, FIFO_DEV_not_dout_2n1s3, 
         FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_0_, 
         FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_1_, 
         FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_2_, 
         FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_3_, 
         FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_4_, 
         FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_5_, 
         FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_6_, 
         FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_7_, nx4093z3, nx4093z2, 
         nx4093z1, nx12521z3, nx11524z1, nx10527z1, nx9530z1, nx8533z1, nx7536z1, 
         nx6539z1, nx5542z1, b_0_, nx37688z1, sclear_and_0_dup_147, 
         sclear_and_1_dup_148, sclear_and_2_dup_149, sclear_and_3_dup_150, 
         sclear_and_4_dup_151, sclear_and_5_dup_152, sclear_and_6_dup_153, 
         sclear_and_7_dup_154, sclear_and_8_dup_155, sclear_and_9_dup_156, 
         sclear_and_10_dup_157, sclear_and_11_dup_158, nx34195z2, nx34318z2, 
         nx27756z1, nx61539z3, nx61539z4, nx61539z2, nx54095z1, nx61539z1, 
         nx34195z1, nx8464z1, nx34318z1, inc_d_3_, inc_d_5_, inc_d_9_, 
         sclear_and_0_dup_719, sclear_and_1_dup_720, sclear_and_2_dup_721, 
         sclear_and_3_dup_722, sclear_and_4_dup_723, sclear_and_5_dup_724, 
         sclear_and_6_dup_725, sclear_and_7_dup_726, sclear_and_8_dup_727, 
         sclear_and_9_dup_728, sclear_and_10_dup_729, sclear_and_11_dup_730, 
         sclear_and_12_dup_731, sclear_and_13_dup_732, sclear_and_14_dup_733, 
         sclear_and_15_dup_734, sclear_and_16_dup_735, sclear_and_17_dup_736, 
         sclear_and_18_dup_737, sclear_and_19_dup_738, sclear_and_20_dup_739, 
         sclear_and_21_dup_740, sclear_and_22_dup_741, sclear_and_23_dup_742, 
         sclear_and_24_dup_743, sclear_and_25_dup_744, sclear_and_26_dup_745, 
         sclear_and_27_dup_746, sclear_and_28_dup_747, sclear_and_29_dup_748, 
         sclear_and_30_dup_749, sclear_and_31_dup_750, sclear_and_32_dup_751, 
         sclear_and_33_dup_752, sclear_and_34_dup_753, sclear_and_35_dup_754, 
         sclear_and_36_dup_755, sclear_and_37_dup_756, sclear_and_38_dup_757, 
         sclear_and_39_dup_758, sclear_and_40_dup_759, sclear_and_41_dup_760, 
         sclear_and_42_dup_761, sclear_and_43_dup_762, sclear_and_44_dup_763, 
         sclear_and_45_dup_764, sclear_and_46_dup_765, sclear_and_47_dup_766, 
         sclear_and_48_dup_767, sclear_and_49_dup_768, sclear_and_50_dup_769, 
         sclear_and_51_dup_770, sclear_and_52_dup_771, sclear_and_53_dup_772, 
         sclear_and_54_dup_773, sclear_and_55_dup_774, sclear_and_56_dup_775, 
         sclear_and_57_dup_776, sclear_and_58_dup_777, sclear_and_59_dup_778, 
         sclear_and_60_dup_779, sclear_and_61_dup_780, sclear_and_62_dup_781, 
         sclear_and_63_dup_782, nx26032z1, nx16750z1, nx8414z3, NOT_a_10_, 
         nx8414z4, nx11298z2, nx11298z3, nx8414z6, nx49501z4, nx56070z3, 
         nx49501z7, nx34946z4, nx49501z9, nx8414z9, nx8409z4, nx8414z11, 
         nx11504z5, nx7417z3, nx11504z7, nx35506z6, nx11504z13, nx55510z4, 
         nx11504z15, nx40554z3, nx41545z2, nx20284z5, nx41545z4, nx19772z4, 
         nx7423z1, nx7418z1, nx9408z1, nx8415z1, NOT_a_4__dup_3628, NOT_a_4_, 
         NOT_a_4__dup_3622, nx6004z1, nx36778z1, nx31484z2, NOT_a_9_, nx8414z5, 
         nx5753z3, nx36042z2, nx49501z3, nx56070z2, nx32220z2, nx10562z3, 
         nx49501z6, nx34946z3, nx7836z3, nx14918z4, nx49501z8, nx8414z8, 
         nx3006z4, nx19748z3, nx8409z3, nx8414z10, nx9406z2, nx9411z2, nx11504z4, 
         nx7417z2, nx32078z2, nx6418z3, nx11504z6, nx35506z5, nx52784z5, 
         nx55534z4, nx11504z12, nx55510z3, nx52808z3, nx35482z3, nx11504z14, 
         nx40554z2, nx39562z2, nx39557z2, nx41545z1, nx20284z4, nx22498z4, 
         nx65280z3, nx41545z3, nx19772z3, nx42542z1, nx60450z3, 
         NOT_a_3__dup_3640, NOT_a_3__dup_3645, NOT_a_3__dup_3650, 
         NOT_a_3__dup_3655, NOT_a_3__dup_3629, NOT_a_3__dup_3635, NOT_a_3_, 
         NOT_a_3__dup_3623, nx51512z1, nx56806z1, nx31484z1, nx11298z1, nx8414z2, 
         nx5753z2, nx10562z2, nx34946z2, nx7836z2, nx14918z3, nx49501z5, 
         nx39776z3, nx3006z3, nx8409z2, nx7411z1, nx7417z1, nx32078z1, nx6418z2, 
         nx11504z3, nx35506z4, nx52784z4, nx55534z3, nx41557z1, nx11504z11, 
         nx40554z1, nx39562z1, nx39557z1, nx20284z3, nx22498z3, nx65280z2, 
         NOT_a_2__dup_3641, NOT_a_2__dup_3646, NOT_a_2__dup_3651, 
         NOT_a_2__dup_3656, NOT_a_2__dup_3630, NOT_a_2__dup_3636, NOT_a_2_, 
         NOT_a_2__dup_3624, nx8414z1, nx5753z1, nx36042z1, nx52248z1, nx56070z1, 
         nx32220z1, nx10562z1, nx12192z1, nx35506z2, nx52784z2, nx14918z2, 
         nx49501z2, nx39776z2, nx3006z2, nx19748z2, nx8409z1, nx8414z7, nx9406z1, 
         nx9411z1, nx2470z2, nx6418z1, NOT_a_7_, nx35506z3, nx52784z3, nx55534z2, 
         nx32756z2, nx55510z2, nx52808z2, nx35482z2, NOT_a_1__dup_3642, 
         NOT_a_1__dup_3647, NOT_a_1__dup_3652, NOT_a_1__dup_3657, 
         NOT_a_1__dup_3631, NOT_a_1__dup_3637, NOT_a_1_, NOT_a_1__dup_3625, 
         nx19772z2, nx46881z2, nx60450z2, nx27840z2, nx14942z2, nx7812z2, 
         nx34970z2, nx34946z1, nx7836z1, nx14918z1, nx49501z1, nx39776z1, 
         nx3006z1, nx19748z1, NOT_a_0__dup_3643, NOT_a_0__dup_3648, 
         NOT_a_0__dup_3653, NOT_a_0__dup_3658, NOT_a_0__dup_3632, 
         NOT_a_0__dup_3638, NOT_a_0_, NOT_a_0__dup_3626, nx7276z1, nx20284z2, 
         nx22498z2, nx23010z2, nx35506z1, nx52784z1, nx55534z1, nx32756z1, 
         nx55510z1, nx52808z1, nx35482z1, nx28937z1, nx60340z1, nx47978z1, 
         nx40312z1, nx2470z1, nx20284z1, nx22498z1, nx65280z1, nx23010z1, 
         nx19772z1, nx46881z1, nx60450z1, nx27840z1, nx14942z1, nx7812z1, 
         nx34970z1, nx12216z1, nx10538z1, nx32244z1, nx56046z1, nx8373z1, 
         nx15368z1, nx27414z1, nx60876z1, sclear_and_0_dup_114, 
         sclear_and_1_dup_115, sclear_and_2_dup_116, sclear_and_3_dup_117, 
         sclear_and_4_dup_118, sclear_and_5_dup_119, sclear_and_6_dup_120, 
         sclear_and_7_dup_121, sclear_and_8_dup_122, nx52196z2, nx24762z1, 
         nx18020z1, nx38048z1, nx52196z1, nx57089z1, nx31201z1, 
         inc_d_3__dup_2781, inc_d_5__dup_2783, inc_d_8__dup_2786, nx32158z1, 
         inc_d_0__dup_2797, inc_d_1__dup_2798, inc_d_2__dup_2799, 
         inc_d_3__dup_2800, inc_d_4__dup_2801, inc_d_5__dup_2802, 
         inc_d_6__dup_2803, inc_d_7__dup_2804, nx54164z2, nx50324z3, nx57994z3, 
         a_0__dup_274, nx47598z1, a_0__dup_276, nx27570z1, nx50324z1, nx57994z1, 
         nx50324z2, a_0__dup_2819, nx54164z1, nx57994z2, incdec_mux_1_dup_99, 
         incdec_mux_2_dup_100, incdec_mux_3_dup_101, incdec_mux_4_dup_102, 
         incdec_mux_5_dup_103, incdec_mux_6_dup_104, incdec_mux_7_dup_105, 
         nx23410z1, nx3438z4, nx10507z2, nx9510z10, nx9510z2, nx9510z8, 
         nx36622z2, nx3438z2, nx18636z2, nx45632z1, nx44635z1, nx43638z1, 
         nx42641z1, nx41644z1, nx40647z1, nx39650z1, nx43638z2, nx40647z3, 
         nx39650z3, nx40647z2, nx39650z2, nx15492z4, nx59980z1, nx37353z2, 
         nx19403z2, nx2452z2, nx19403z3, nx50038z2, nx45412z2, nx63362z2, 
         nx15776z2, nx63362z3, nx32727z2, nx50677z2, nx2092z2, nx9565z2, 
         nx2092z3, nx27515z2, nx37353z3, nx44466z2, nx62416z3, nx62416z2, 
         nx13831z3, nx13831z2, nx37353z4, nx36356z2, nx35359z2, nx49948z1, 
         nx34362z2, nx33365z2, nx32368z2, nx30372z2, nx32368z3, nx29375z2, 
         nx28378z2, nx27381z2, nx26384z2, nx27381z3, nx25387z2, nx33365z3, 
         nx24390z2, nx23393z3, nx23393z2, nx22396z3, nx22396z2, nx21399z3, 
         nx21399z2, nx31781z3, nx31781z2, nx35840z1, nx36837z1, nx36837z2, 
         nx37834z1, nx37834z2, nx38831z1, nx38831z2, nx39828z1, nx39828z2, 
         nx40825z1, nx40825z2, nx41822z1, nx41822z2, nx42819z1, nx43816z1, 
         nx43816z2, nx44813z1, nx44813z2, nx32187z1, nx32187z2, nx31190z1, 
         nx31190z2, nx30193z1, nx30193z2, nx29196z1, nx29196z2, nx28199z1, 
         nx28199z2, nx27202z1, nx27202z2, nx26205z1, nx26205z2, nx25208z1, 
         nx25208z2, nx24211z1, nx24211z2, nx23214z1, nx23214z2, nx21218z1, 
         nx21218z2, nx20221z1, nx20221z2, nx19224z1, nx19224z2, nx18227z1, 
         nx18227z2, nx17230z1, nx17230z2, nx16233z1, nx16233z2, nx15236z1, 
         nx15236z2, nx14239z1, nx14239z2, nx13242z1, nx13242z2, nx12245z1, 
         nx12245z2, nx10249z1, nx10249z2, nx9252z1, nx9252z2, nx8255z1, nx8255z2, 
         nx7258z1, nx7258z2, nx6261z1, nx6261z2, nx5264z1, nx5264z2, nx4267z1, 
         nx4267z2, nx3270z1, nx3270z2, nx2273z1, nx2273z2, nx1276z1, nx1276z2, 
         nx64816z1, nx64816z2, nx63819z1, nx63819z2, nx62822z1, nx62822z2, 
         nx61825z1, nx61825z2, nx60828z1, nx60828z2, nx59831z1, nx59831z2, 
         nx58834z1, nx58834z2, nx57837z1, nx57837z2, nx56840z1, nx56840z2, 
         nx55843z1, nx55843z2, nx53847z1, nx53847z2, nx52850z1, nx52850z2, 
         nx51853z1, nx51853z2, nx50856z1, nx50856z2, nx49859z1, nx49859z2, 
         nx48862z1, nx48862z2, nx47865z1, nx47865z2, nx46868z1, nx46868z2, 
         nx45871z1, nx45871z2, nx44874z1, nx44874z2, nx42878z1, nx42878z2, 
         nx41881z1, nx41881z2, nx40884z1, nx40884z2, nx39887z1, nx39887z2, 
         nx38890z1, nx38890z2, nx37893z1, nx37893z2, nx36896z1, nx36896z2, 
         nx35899z1, nx35899z2, nx34902z1, nx34902z2, nx33905z1, nx33905z2, 
         nx31909z1, nx31909z2, nx30912z1, nx30912z2, nx29915z1, nx29915z2, 
         nx28918z1, nx28918z2, nx27921z1, nx27921z2, nx26924z1, nx26924z2, 
         nx25927z1, nx25927z2, nx24930z1, nx24930z2, nx23933z1, nx22936z1, 
         nx20940z1, nx19943z1, nx18946z1, nx17949z1, nx16952z1, nx15955z1, 
         nx14958z1, nx13961z1, nx12964z1, nx11967z1, nx9971z1, nx8974z1, 
         nx7977z1, nx58629z1, nx59626z1, nx60623z1, nx61620z1, nx21254z1, 
         nx20257z1, nx19260z1, nx18263z1, nx17266z1, nx16269z1, nx15272z1, 
         nx14275z1, nx13278z1, nx12281z1, nx4121z1, nx3124z1, nx2127z1, nx1130z1, 
         nx133z1, nx64672z1, nx63675z1, nx62678z1, nx61681z1, nx60684z1, 
         nx58688z1, nx57691z1, nx56694z1, nx55697z1, nx54700z1, nx53703z1, 
         nx52706z1, nx51709z1, nx50712z1, nx49715z1, nx47719z1, nx46722z1, 
         nx45725z1, nx44728z1, nx43731z1, nx42734z1, nx41737z1, nx40740z1, 
         nx39743z1, nx38746z1, nx36750z1, nx35753z1, nx34756z1, nx33759z1, 
         nx32762z1, nx31765z1, nx30768z1, nx29771z1, nx28774z1, nx27777z1, 
         nx25781z1, nx24784z1, nx23787z1, nx22790z1, nx21793z1, nx20796z1, 
         nx19799z1, nx18802z1, nx17805z1, nx16808z2, nx14812z1, nx13815z1, 
         nx12818z1, nx11821z1, nx10824z1, nx9827z1, nx8830z1, nx7833z1, nx6836z1, 
         nx5839z1, nx3843z1, nx2846z1, nx1849z1, nx852z1, nx65391z1, nx64394z1, 
         nx63397z1, nx62400z1, nx61403z1, nx60406z1, nx58410z1, nx57413z1, 
         nx56416z1, nx55419z1, nx54422z1, nx53425z1, nx52428z1, nx51431z1, 
         nx50434z1, nx49437z1, nx47441z1, nx46444z1, nx45447z1, nx44450z1, 
         nx43453z1, nx42456z1, nx41459z1, nx40462z1, nx39465z1, nx38468z1, 
         nx27151z1, nx28148z1, nx29145z1, nx30142z1, nx31139z1, nx32136z1, 
         nx33133z1, nx34130z1, nx24478z1, nx23481z1, nx21487z1, nx20490z1, 
         nx19493z1, nx18496z1, nx16502z1, nx48379z1, nx49376z1, nx52367z1, 
         nx53364z1, nx56355z1, nx58351z1, nx59348z1, nx61342z1, nx62339z1, 
         nx63336z1, nx64333z1, nx65330z1, nx4781z1, nx5778z1, nx6775z1, nx8769z1, 
         nx10763z1, nx14753z1, nx17744z1, nx19738z1, nx21732z1, nx25722z1, 
         nx28713z1, nx30707z1, nx32701z1, nx33698z1, nx34695z1, nx39682z1, 
         nx40679z1, nx43670z1, nx44667z1, nx45664z1, nx47660z1, nx49654z1, 
         nx52645z1, nx53642z1, nx54639z1, NOT_a_2__dup_4701, NOT_a_1__dup_4702, 
         nx12216z2, nx15492z6, nx15492z7, nx15492z8, nx9510z5, nx9510z4, 
         nx9510z7, nx9510z6, nx11504z9, nx11504z8, nx10507z4, nx11504z17, 
         nx11504z16, nx11504z10, nx11504z2, nx11504z20, nx11504z21, nx11504z19, 
         nx41852z2, nx41852z1, nx41852z3, nx41852z4, nx54297z2, nx54297z1, 
         nx54297z3, nx54297z4, nx48026z2, nx48026z1, nx48026z3, nx47029z2, 
         nx47029z1, nx47029z3, nx46032z2, nx46032z1, nx46032z3, nx45035z2, 
         nx45035z1, nx45035z3, nx44038z2, nx44038z1, nx44038z3, nx43041z2, 
         nx43041z1, nx43041z3, nx42044z2, nx42044z1, nx42044z3, nx41047z2, 
         nx41047z1, nx41047z3, nx27414z3, nx27414z2, nx60876z3, nx60876z2, 
         nx8373z2, nx15368z2, nx15368z3, nx10538z2, nx32244z2, nx56046z2, 
         nx7969z1, nx19668z1, nx55223z1, ENCR_DEV_rtlc15_PS14_n166, nx37353z1, 
         nx36356z1, nx35359z1, nx34362z1, nx33365z1, nx32368z1, nx30372z1, 
         nx29375z1, nx28378z1, nx27381z1, nx26384z1, nx25387z1, nx24390z1, 
         nx23393z1, nx22396z1, nx21399z1, nx19403z1, nx18406z1, nx17409z1, 
         nx16412z1, nx15415z1, nx14418z1, nx13421z1, nx12424z1, nx11427z1, 
         nx10430z1, nx8434z1, nx7437z1, nx6440z1, nx5443z1, nx4446z1, nx3449z1, 
         nx2452z1, nx1455z1, nx458z1, nx64997z1, nx63001z1, nx62004z1, nx61007z1, 
         nx60010z1, nx59013z1, nx58016z1, nx57019z1, nx56022z1, nx55025z1, 
         nx54028z1, nx52032z1, nx51035z1, nx50038z1, nx49041z1, nx48044z1, 
         nx47047z1, nx46050z1, nx45053z1, nx44056z1, nx43059z1, nx37436z1, 
         nx38433z1, nx39430z1, nx40427z1, nx41424z1, nx42421z1, nx43418z1, 
         nx44415z1, nx45412z1, nx46409z1, nx48405z1, nx49402z1, nx50399z1, 
         nx51396z1, nx52393z1, nx53390z1, nx54387z1, nx55384z1, nx56381z1, 
         nx57378z1, nx59374z1, nx60371z1, nx61368z1, nx62365z1, nx63362z1, 
         nx64359z1, nx65356z1, nx817z1, nx1814z1, nx2811z1, nx4807z1, nx5804z1, 
         nx6801z1, nx7798z1, nx8795z1, nx9792z1, nx10789z1, nx11786z1, nx12783z1, 
         nx13780z1, nx15776z1, nx16773z1, nx17770z1, nx18767z1, nx19764z1, 
         nx20761z1, nx21758z1, nx22755z1, nx23752z1, nx24749z1, nx26745z1, 
         nx27742z1, nx28739z1, nx29736z1, nx30733z1, nx31730z1, nx32727z1, 
         nx33724z1, nx34721z1, nx35718z1, nx37714z1, nx38711z1, nx39708z1, 
         nx40705z1, nx41702z1, nx42699z1, nx43696z1, nx44693z1, nx45690z1, 
         nx46687z1, nx48683z1, nx49680z1, nx50677z1, nx51674z1, nx52671z1, 
         nx53668z1, nx54665z1, nx55662z1, nx56659z1, nx57656z1, nx59652z1, 
         nx60649z1, nx61646z1, nx62643z1, nx63640z1, nx64637z1, nx98z1, nx1095z1, 
         nx2092z1, nx3089z1, nx5085z1, nx6082z1, nx7079z1, nx8076z1, nx9073z1, 
         nx10070z1, nx11067z1, nx12064z1, nx13061z1, nx14058z1, nx5577z1, 
         nx6574z1, nx7571z1, nx8568z1, nx9565z1, nx10562z4, nx11559z1, nx12556z1, 
         nx13553z1, nx14550z1, nx16546z1, nx17543z1, nx18540z1, nx19537z1, 
         nx20534z1, nx21531z1, nx22528z1, nx23525z1, nx24522z1, nx25519z1, 
         nx27515z1, nx28512z1, nx29509z1, nx30506z1, nx31503z1, nx32500z1, 
         nx33497z1, nx34494z1, nx35491z1, nx36488z1, nx38484z1, nx39481z1, 
         nx40478z1, nx41475z1, nx42472z1, nx43469z1, nx44466z1, nx45463z1, 
         nx46460z1, nx47457z1, nx49453z1, nx50450z1, nx51447z1, nx52444z1, 
         nx53441z1, nx54438z1, nx55435z1, nx56432z1, nx57429z1, nx58426z1, 
         nx60422z1, nx61419z1, nx62416z1, nx63413z1, nx64410z1, nx65407z1, 
         nx868z1, nx1865z1, nx2862z1, nx3859z1, nx5855z1, nx6852z1, nx7849z1, 
         nx8846z1, nx9843z1, nx10840z1, nx11837z1, nx12834z1, nx13831z1, 
         nx14828z1, nx16824z1, nx17821z1, nx18818z1, nx19815z1, nx20812z1, 
         nx21809z1, nx22806z1, nx23803z1, nx24800z1, nx25797z1, nx27793z1, 
         nx28790z1, nx29787z1, nx30784z1, nx31781z1, nx32778z1, nx33775z1, 
         nx34772z1, nx35769z1, nx36766z1, nx48358z1, nx47361z1, nx46364z1, 
         nx45367z1, nx44370z1, nx43373z1, nx42376z1, nx41379z1, nx40382z1, 
         nx39385z1, nx12521z2, FIFO_DEV_rtlc14_X_0_n123, nx45632z2, nx22484z1, 
         nx25475z1, nx5542z3, nx6539z3, nx7536z3, nx8533z3, nx9530z3, nx10527z3, 
         nx11524z3, nx12521z7, nx35840z2, nx42819z2, nx25475z3, nx22484z3, 
         nx17499z1, nx17499z2, nx47382z1, nx47382z2, nx50373z1, nx50373z2, 
         nx51370z1, nx51370z2, nx54361z1, nx54361z2, nx55358z1, nx55358z2, 
         nx60345z1, nx60345z2, nx791z1, nx791z2, nx1788z1, nx1788z2, nx3784z1, 
         nx3784z2, nx7772z1, nx7772z2, nx9766z1, nx9766z2, nx11760z1, nx11760z2, 
         nx12757z1, nx12757z2, nx15750z1, nx15750z2, nx16747z1, nx16747z2, 
         nx18741z1, nx18741z2, nx20735z1, nx20735z2, nx22729z1, nx22729z2, 
         nx23726z1, nx23726z2, nx26719z1, nx26719z2, nx27716z1, nx27716z2, 
         nx29710z1, nx29710z2, nx31704z1, nx31704z2, nx36691z1, nx36691z2, 
         nx37688z2, nx37688z3, nx38685z1, nx38685z2, nx41676z1, nx41676z2, 
         nx42673z1, nx42673z2, nx48657z1, nx48657z2, nx50651z1, nx50651z2, 
         nx51648z1, nx51648z2, nx55636z1, nx55636z2, nx56633z1, nx56633z2, 
         nx35127z1, nx35127z2, nx36124z1, nx36124z2, nx38120z1, nx38120z2, 
         nx11504z18, nx65298z1, nx16808z1, nx32158z3, nx12521z9, nx12521z10, 
         ENCR_DEV_prev_6__int, NOT_FIFO_DEV_rtlc5n43_int, b_0__int, 
         NOT_ENCR_DEV_rtlcn261_int, NOT_ENCR_DEV_rtlc12n435__repl0, 
         NOT_ENCR_DEV_rtlc12n435__repl1, NOT_ENCR_DEV_rtlc12n435__repl2, 
         FIFO_DEV_rtlc_radd_N1_5___repl0, FIFO_DEV_rtlc_radd_N1_5___repl1, 
         FIFO_DEV_rtlc_radd_N1_3___repl0, FIFO_DEV_rtlc_radd_N1_2___repl0, 
         FIFO_DEV_rtlc_radd_N1_2___repl1, FIFO_DEV_rtlc_radd_N1_2___repl2, 
         FIFO_DEV_rtlc_radd_N1_1___repl0, FIFO_DEV_rtlc_radd_N1_0___repl0, 
         NOT_ENCR_DEV_rtlc15n971__repl0, NOT_ENCR_DEV_rtlc15n971__repl1, 
         NOT_ENCR_DEV_rtlc15n971__repl2, NOT_ENCR_DEV_rtlc15n971__repl3, 
         NOT_ENCR_DEV_rtlc15n971__repl4, NOT_ENCR_DEV_rtlc15n971__repl5, 
         ENCR_DEV_prev_5___repl0, ENCR_DEV_prev_5___repl1, 
         ENCR_DEV_prev_5___repl2, NOT_ENCR_DEV_rtlc15n968__repl0, 
         NOT_ENCR_DEV_rtlc15n968__repl1, NOT_ENCR_DEV_rtlc15n968__repl2, 
         NOT_ENCR_DEV_rtlc15n968__repl3, NOT_ENCR_DEV_rtlc15n968__repl4, 
         ENCR_DEV_prev_1___repl0, ENCR_DEV_prev_1___repl1, 
         ENCR_DEV_prev_1___repl2, ENCR_DEV_prev_1___repl3, 
         ENCR_DEV_prev_1___repl4, ENCR_DEV_rtlcn483__repl0, 
         ENCR_DEV_rtlcn483__repl1, ENCR_DEV_rtlcn483__repl2, 
         ENCR_DEV_prev_8___repl0, ENCR_DEV_prev_8___repl1, 
         ENCR_DEV_prev_8___repl2, ENCR_DEV_prev_8___repl3, 
         ENCR_DEV_prev_8___repl4, ENCR_DEV_prev_8___repl5, 
         ENCR_DEV_prev_8___repl6;
    wire [279:0] \$dummy ;




    mux_256_0 FIFO_DEV_dout_mux_2i1 (.a ({FIFO_DEV_rtlc_msr_n3[255],
              FIFO_DEV_rtlc_msr_n3[254],FIFO_DEV_rtlc_msr_n3[253],
              FIFO_DEV_rtlc_msr_n3[252],FIFO_DEV_rtlc_msr_n3[251],
              FIFO_DEV_rtlc_msr_n3[250],FIFO_DEV_rtlc_msr_n3[249],
              FIFO_DEV_rtlc_msr_n3[248],FIFO_DEV_rtlc_msr_n3[247],
              FIFO_DEV_rtlc_msr_n3[246],FIFO_DEV_rtlc_msr_n3[245],
              FIFO_DEV_rtlc_msr_n3[244],FIFO_DEV_rtlc_msr_n3[243],
              FIFO_DEV_rtlc_msr_n3[242],FIFO_DEV_rtlc_msr_n3[241],
              FIFO_DEV_rtlc_msr_n3[240],FIFO_DEV_rtlc_msr_n3[239],
              FIFO_DEV_rtlc_msr_n3[238],FIFO_DEV_rtlc_msr_n3[237],
              FIFO_DEV_rtlc_msr_n3[236],FIFO_DEV_rtlc_msr_n3[235],
              FIFO_DEV_rtlc_msr_n3[234],FIFO_DEV_rtlc_msr_n3[233],
              FIFO_DEV_rtlc_msr_n3[232],FIFO_DEV_rtlc_msr_n3[231],
              FIFO_DEV_rtlc_msr_n3[230],FIFO_DEV_rtlc_msr_n3[229],
              FIFO_DEV_rtlc_msr_n3[228],FIFO_DEV_rtlc_msr_n3[227],
              FIFO_DEV_rtlc_msr_n3[226],FIFO_DEV_rtlc_msr_n3[225],
              FIFO_DEV_rtlc_msr_n3[224],FIFO_DEV_rtlc_msr_n3[223],
              FIFO_DEV_rtlc_msr_n3[222],FIFO_DEV_rtlc_msr_n3[221],
              FIFO_DEV_rtlc_msr_n3[220],FIFO_DEV_rtlc_msr_n3[219],
              FIFO_DEV_rtlc_msr_n3[218],FIFO_DEV_rtlc_msr_n3[217],
              FIFO_DEV_rtlc_msr_n3[216],FIFO_DEV_rtlc_msr_n3[215],
              FIFO_DEV_rtlc_msr_n3[214],FIFO_DEV_rtlc_msr_n3[213],
              FIFO_DEV_rtlc_msr_n3[212],FIFO_DEV_rtlc_msr_n3[211],
              FIFO_DEV_rtlc_msr_n3[210],FIFO_DEV_rtlc_msr_n3[209],
              FIFO_DEV_rtlc_msr_n3[208],FIFO_DEV_rtlc_msr_n3[207],
              FIFO_DEV_rtlc_msr_n3[206],FIFO_DEV_rtlc_msr_n3[205],
              FIFO_DEV_rtlc_msr_n3[204],FIFO_DEV_rtlc_msr_n3[203],
              FIFO_DEV_rtlc_msr_n3[202],FIFO_DEV_rtlc_msr_n3[201],
              FIFO_DEV_rtlc_msr_n3[200],FIFO_DEV_rtlc_msr_n3[199],
              FIFO_DEV_rtlc_msr_n3[198],FIFO_DEV_rtlc_msr_n3[197],
              FIFO_DEV_rtlc_msr_n3[196],FIFO_DEV_rtlc_msr_n3[195],
              FIFO_DEV_rtlc_msr_n3[194],FIFO_DEV_rtlc_msr_n3[193],
              FIFO_DEV_rtlc_msr_n3[192],FIFO_DEV_rtlc_msr_n3[191],
              FIFO_DEV_rtlc_msr_n3[190],FIFO_DEV_rtlc_msr_n3[189],
              FIFO_DEV_rtlc_msr_n3[188],FIFO_DEV_rtlc_msr_n3[187],
              FIFO_DEV_rtlc_msr_n3[186],FIFO_DEV_rtlc_msr_n3[185],
              FIFO_DEV_rtlc_msr_n3[184],FIFO_DEV_rtlc_msr_n3[183],
              FIFO_DEV_rtlc_msr_n3[182],FIFO_DEV_rtlc_msr_n3[181],
              FIFO_DEV_rtlc_msr_n3[180],FIFO_DEV_rtlc_msr_n3[179],
              FIFO_DEV_rtlc_msr_n3[178],FIFO_DEV_rtlc_msr_n3[177],
              FIFO_DEV_rtlc_msr_n3[176],FIFO_DEV_rtlc_msr_n3[175],
              FIFO_DEV_rtlc_msr_n3[174],FIFO_DEV_rtlc_msr_n3[173],
              FIFO_DEV_rtlc_msr_n3[172],FIFO_DEV_rtlc_msr_n3[171],
              FIFO_DEV_rtlc_msr_n3[170],FIFO_DEV_rtlc_msr_n3[169],
              FIFO_DEV_rtlc_msr_n3[168],FIFO_DEV_rtlc_msr_n3[167],
              FIFO_DEV_rtlc_msr_n3[166],FIFO_DEV_rtlc_msr_n3[165],
              FIFO_DEV_rtlc_msr_n3[164],FIFO_DEV_rtlc_msr_n3[163],
              FIFO_DEV_rtlc_msr_n3[162],FIFO_DEV_rtlc_msr_n3[161],
              FIFO_DEV_rtlc_msr_n3[160],FIFO_DEV_rtlc_msr_n3[159],
              FIFO_DEV_rtlc_msr_n3[158],FIFO_DEV_rtlc_msr_n3[157],
              FIFO_DEV_rtlc_msr_n3[156],FIFO_DEV_rtlc_msr_n3[155],
              FIFO_DEV_rtlc_msr_n3[154],FIFO_DEV_rtlc_msr_n3[153],
              FIFO_DEV_rtlc_msr_n3[152],FIFO_DEV_rtlc_msr_n3[151],
              FIFO_DEV_rtlc_msr_n3[150],FIFO_DEV_rtlc_msr_n3[149],
              FIFO_DEV_rtlc_msr_n3[148],FIFO_DEV_rtlc_msr_n3[147],
              FIFO_DEV_rtlc_msr_n3[146],FIFO_DEV_rtlc_msr_n3[145],
              FIFO_DEV_rtlc_msr_n3[144],FIFO_DEV_rtlc_msr_n3[143],
              FIFO_DEV_rtlc_msr_n3[142],FIFO_DEV_rtlc_msr_n3[141],
              FIFO_DEV_rtlc_msr_n3[140],FIFO_DEV_rtlc_msr_n3[139],
              FIFO_DEV_rtlc_msr_n3[138],FIFO_DEV_rtlc_msr_n3[137],
              FIFO_DEV_rtlc_msr_n3[136],FIFO_DEV_rtlc_msr_n3[135],
              FIFO_DEV_rtlc_msr_n3[134],FIFO_DEV_rtlc_msr_n3[133],
              FIFO_DEV_rtlc_msr_n3[132],FIFO_DEV_rtlc_msr_n3[131],
              FIFO_DEV_rtlc_msr_n3[130],FIFO_DEV_rtlc_msr_n3[129],
              FIFO_DEV_rtlc_msr_n3[128],FIFO_DEV_rtlc_msr_n3[127],
              FIFO_DEV_rtlc_msr_n3[126],FIFO_DEV_rtlc_msr_n3[125],
              FIFO_DEV_rtlc_msr_n3[124],FIFO_DEV_rtlc_msr_n3[123],
              FIFO_DEV_rtlc_msr_n3[122],FIFO_DEV_rtlc_msr_n3[121],
              FIFO_DEV_rtlc_msr_n3[120],FIFO_DEV_rtlc_msr_n3[119],
              FIFO_DEV_rtlc_msr_n3[118],FIFO_DEV_rtlc_msr_n3[117],
              FIFO_DEV_rtlc_msr_n3[116],FIFO_DEV_rtlc_msr_n3[115],
              FIFO_DEV_rtlc_msr_n3[114],FIFO_DEV_rtlc_msr_n3[113],
              FIFO_DEV_rtlc_msr_n3[112],FIFO_DEV_rtlc_msr_n3[111],
              FIFO_DEV_rtlc_msr_n3[110],FIFO_DEV_rtlc_msr_n3[109],
              FIFO_DEV_rtlc_msr_n3[108],FIFO_DEV_rtlc_msr_n3[107],
              FIFO_DEV_rtlc_msr_n3[106],FIFO_DEV_rtlc_msr_n3[105],
              FIFO_DEV_rtlc_msr_n3[104],FIFO_DEV_rtlc_msr_n3[103],
              FIFO_DEV_rtlc_msr_n3[102],FIFO_DEV_rtlc_msr_n3[101],
              FIFO_DEV_rtlc_msr_n3[100],FIFO_DEV_rtlc_msr_n3[99],
              FIFO_DEV_rtlc_msr_n3[98],FIFO_DEV_rtlc_msr_n3[97],
              FIFO_DEV_rtlc_msr_n3[96],FIFO_DEV_rtlc_msr_n3[95],
              FIFO_DEV_rtlc_msr_n3[94],FIFO_DEV_rtlc_msr_n3[93],
              FIFO_DEV_rtlc_msr_n3[92],FIFO_DEV_rtlc_msr_n3[91],
              FIFO_DEV_rtlc_msr_n3[90],FIFO_DEV_rtlc_msr_n3[89],
              FIFO_DEV_rtlc_msr_n3[88],FIFO_DEV_rtlc_msr_n3[87],
              FIFO_DEV_rtlc_msr_n3[86],FIFO_DEV_rtlc_msr_n3[85],
              FIFO_DEV_rtlc_msr_n3[84],FIFO_DEV_rtlc_msr_n3[83],
              FIFO_DEV_rtlc_msr_n3[82],FIFO_DEV_rtlc_msr_n3[81],
              FIFO_DEV_rtlc_msr_n3[80],FIFO_DEV_rtlc_msr_n3[79],
              FIFO_DEV_rtlc_msr_n3[78],FIFO_DEV_rtlc_msr_n3[77],
              FIFO_DEV_rtlc_msr_n3[76],FIFO_DEV_rtlc_msr_n3[75],
              FIFO_DEV_rtlc_msr_n3[74],FIFO_DEV_rtlc_msr_n3[73],
              FIFO_DEV_rtlc_msr_n3[72],FIFO_DEV_rtlc_msr_n3[71],
              FIFO_DEV_rtlc_msr_n3[70],FIFO_DEV_rtlc_msr_n3[69],
              FIFO_DEV_rtlc_msr_n3[68],FIFO_DEV_rtlc_msr_n3[67],
              FIFO_DEV_rtlc_msr_n3[66],FIFO_DEV_rtlc_msr_n3[65],
              FIFO_DEV_rtlc_msr_n3[64],FIFO_DEV_rtlc_msr_n3[63],
              FIFO_DEV_rtlc_msr_n3[62],FIFO_DEV_rtlc_msr_n3[61],
              FIFO_DEV_rtlc_msr_n3[60],FIFO_DEV_rtlc_msr_n3[59],
              FIFO_DEV_rtlc_msr_n3[58],FIFO_DEV_rtlc_msr_n3[57],
              FIFO_DEV_rtlc_msr_n3[56],FIFO_DEV_rtlc_msr_n3[55],
              FIFO_DEV_rtlc_msr_n3[54],FIFO_DEV_rtlc_msr_n3[53],
              FIFO_DEV_rtlc_msr_n3[52],FIFO_DEV_rtlc_msr_n3[51],
              FIFO_DEV_rtlc_msr_n3[50],FIFO_DEV_rtlc_msr_n3[49],
              FIFO_DEV_rtlc_msr_n3[48],FIFO_DEV_rtlc_msr_n3[47],
              FIFO_DEV_rtlc_msr_n3[46],FIFO_DEV_rtlc_msr_n3[45],
              FIFO_DEV_rtlc_msr_n3[44],FIFO_DEV_rtlc_msr_n3[43],
              FIFO_DEV_rtlc_msr_n3[42],FIFO_DEV_rtlc_msr_n3[41],
              FIFO_DEV_rtlc_msr_n3[40],FIFO_DEV_rtlc_msr_n3[39],
              FIFO_DEV_rtlc_msr_n3[38],FIFO_DEV_rtlc_msr_n3[37],
              FIFO_DEV_rtlc_msr_n3[36],FIFO_DEV_rtlc_msr_n3[35],
              FIFO_DEV_rtlc_msr_n3[34],FIFO_DEV_rtlc_msr_n3[33],
              FIFO_DEV_rtlc_msr_n3[32],FIFO_DEV_rtlc_msr_n3[31],
              FIFO_DEV_rtlc_msr_n3[30],FIFO_DEV_rtlc_msr_n3[29],
              FIFO_DEV_rtlc_msr_n3[28],FIFO_DEV_rtlc_msr_n3[27],
              FIFO_DEV_rtlc_msr_n3[26],FIFO_DEV_rtlc_msr_n3[25],
              FIFO_DEV_rtlc_msr_n3[24],FIFO_DEV_rtlc_msr_n3[23],
              FIFO_DEV_rtlc_msr_n3[22],FIFO_DEV_rtlc_msr_n3[21],
              FIFO_DEV_rtlc_msr_n3[20],FIFO_DEV_rtlc_msr_n3[19],
              FIFO_DEV_rtlc_msr_n3[18],FIFO_DEV_rtlc_msr_n3[17],
              FIFO_DEV_rtlc_msr_n3[16],FIFO_DEV_rtlc_msr_n3[15],
              FIFO_DEV_rtlc_msr_n3[14],FIFO_DEV_rtlc_msr_n3[13],
              FIFO_DEV_rtlc_msr_n3[12],FIFO_DEV_rtlc_msr_n3[11],
              FIFO_DEV_rtlc_msr_n3[10],FIFO_DEV_rtlc_msr_n3[9],
              FIFO_DEV_rtlc_msr_n3[8],FIFO_DEV_rtlc_msr_n3[7],
              FIFO_DEV_rtlc_msr_n3[6],FIFO_DEV_rtlc_msr_n3[5],
              FIFO_DEV_rtlc_msr_n3[4],FIFO_DEV_rtlc_msr_n3[3],
              FIFO_DEV_rtlc_msr_n3[2],FIFO_DEV_rtlc_msr_n3[1],
              FIFO_DEV_rtlc_msr_n3[0]}), .b ({\$dummy [0],\$dummy [1],
              \$dummy [2],\$dummy [3],\$dummy [4],\$dummy [5],\$dummy [6],
              \$dummy [7],\$dummy [8],\$dummy [9],\$dummy [10],\$dummy [11],
              \$dummy [12],\$dummy [13],\$dummy [14],\$dummy [15],\$dummy [16],
              \$dummy [17],\$dummy [18],\$dummy [19],\$dummy [20],\$dummy [21],
              \$dummy [22],\$dummy [23],\$dummy [24],\$dummy [25],\$dummy [26],
              \$dummy [27],\$dummy [28],\$dummy [29],\$dummy [30],\$dummy [31],
              \$dummy [32],\$dummy [33],\$dummy [34],\$dummy [35],\$dummy [36],
              \$dummy [37],\$dummy [38],\$dummy [39],\$dummy [40],\$dummy [41],
              \$dummy [42],\$dummy [43],\$dummy [44],\$dummy [45],\$dummy [46],
              \$dummy [47],\$dummy [48],\$dummy [49],\$dummy [50],\$dummy [51],
              \$dummy [52],\$dummy [53],\$dummy [54],\$dummy [55],\$dummy [56],
              \$dummy [57],\$dummy [58],\$dummy [59],\$dummy [60],\$dummy [61],
              \$dummy [62],\$dummy [63],\$dummy [64],\$dummy [65],\$dummy [66],
              \$dummy [67],\$dummy [68],\$dummy [69],\$dummy [70],\$dummy [71],
              \$dummy [72],\$dummy [73],\$dummy [74],\$dummy [75],\$dummy [76],
              \$dummy [77],\$dummy [78],\$dummy [79],\$dummy [80],\$dummy [81],
              \$dummy [82],\$dummy [83],\$dummy [84],\$dummy [85],\$dummy [86],
              \$dummy [87],\$dummy [88],\$dummy [89],\$dummy [90],\$dummy [91],
              \$dummy [92],\$dummy [93],\$dummy [94],\$dummy [95],\$dummy [96],
              \$dummy [97],\$dummy [98],\$dummy [99],\$dummy [100],\$dummy [101]
              ,\$dummy [102],\$dummy [103],\$dummy [104],\$dummy [105],
              \$dummy [106],\$dummy [107],\$dummy [108],\$dummy [109],
              \$dummy [110],\$dummy [111],\$dummy [112],\$dummy [113],
              \$dummy [114],\$dummy [115],\$dummy [116],\$dummy [117],
              \$dummy [118],\$dummy [119],\$dummy [120],\$dummy [121],
              \$dummy [122],\$dummy [123],\$dummy [124],\$dummy [125],
              \$dummy [126],\$dummy [127],\$dummy [128],\$dummy [129],
              \$dummy [130],\$dummy [131],\$dummy [132],\$dummy [133],
              \$dummy [134],\$dummy [135],\$dummy [136],\$dummy [137],
              \$dummy [138],\$dummy [139],\$dummy [140],\$dummy [141],
              \$dummy [142],\$dummy [143],\$dummy [144],\$dummy [145],
              \$dummy [146],\$dummy [147],\$dummy [148],\$dummy [149],
              \$dummy [150],\$dummy [151],\$dummy [152],\$dummy [153],
              \$dummy [154],\$dummy [155],\$dummy [156],\$dummy [157],
              \$dummy [158],\$dummy [159],\$dummy [160],\$dummy [161],
              \$dummy [162],\$dummy [163],\$dummy [164],\$dummy [165],
              \$dummy [166],\$dummy [167],\$dummy [168],\$dummy [169],
              \$dummy [170],\$dummy [171],\$dummy [172],\$dummy [173],
              \$dummy [174],\$dummy [175],\$dummy [176],\$dummy [177],
              \$dummy [178],\$dummy [179],\$dummy [180],\$dummy [181],
              \$dummy [182],\$dummy [183],\$dummy [184],\$dummy [185],
              \$dummy [186],\$dummy [187],\$dummy [188],\$dummy [189],
              \$dummy [190],\$dummy [191],\$dummy [192],\$dummy [193],
              \$dummy [194],\$dummy [195],\$dummy [196],\$dummy [197],
              \$dummy [198],\$dummy [199],\$dummy [200],\$dummy [201],
              \$dummy [202],\$dummy [203],\$dummy [204],\$dummy [205],
              \$dummy [206],\$dummy [207],\$dummy [208],\$dummy [209],
              \$dummy [210],\$dummy [211],\$dummy [212],\$dummy [213],
              \$dummy [214],\$dummy [215],\$dummy [216],\$dummy [217],
              \$dummy [218],\$dummy [219],\$dummy [220],\$dummy [221],
              \$dummy [222],\$dummy [223],\$dummy [224],\$dummy [225],
              \$dummy [226],\$dummy [227],\$dummy [228],\$dummy [229],
              \$dummy [230],\$dummy [231],\$dummy [232],\$dummy [233],
              \$dummy [234],\$dummy [235],\$dummy [236],\$dummy [237],
              \$dummy [238],\$dummy [239],\$dummy [240],\$dummy [241],
              \$dummy [242],\$dummy [243],\$dummy [244],\$dummy [245],
              \$dummy [246],\$dummy [247],\$dummy [248],FIFO_DEV_rtlc_radd_N1[6]
              ,FIFO_DEV_rtlc_radd_N1[5],FIFO_DEV_rtlc_radd_N1[4],
              FIFO_DEV_rtlc_radd_N1[3],FIFO_DEV_rtlc_radd_N1[2],
              FIFO_DEV_rtlc_radd_N1[1],FIFO_DEV_rtlc_radd_N1[0]}), .d (
              \$dummy [249]), .px994 (nx12521z9), .px775 (nx12521z10), .p_FIFO_DEV_rtlc_radd_N1_5___repl0 (
              FIFO_DEV_rtlc_radd_N1_5___repl0), .p_FIFO_DEV_rtlc_radd_N1_5___repl1 (
              FIFO_DEV_rtlc_radd_N1_5___repl1), .p_FIFO_DEV_rtlc_radd_N1_3___repl0 (
              FIFO_DEV_rtlc_radd_N1_3___repl0), .p_FIFO_DEV_rtlc_radd_N1_2___repl0 (
              FIFO_DEV_rtlc_radd_N1_2___repl0), .p_FIFO_DEV_rtlc_radd_N1_2___repl1 (
              FIFO_DEV_rtlc_radd_N1_2___repl1), .p_FIFO_DEV_rtlc_radd_N1_2___repl2 (
              FIFO_DEV_rtlc_radd_N1_2___repl2), .p_FIFO_DEV_rtlc_radd_N1_1___repl0 (
              FIFO_DEV_rtlc_radd_N1_1___repl0), .p_FIFO_DEV_rtlc_radd_N1_0___repl0 (
              FIFO_DEV_rtlc_radd_N1_0___repl0)) ;
    ram_dq_8_0 FIFO_DEV_fifomem (.wr_data1 ({STREAM[7],STREAM[6],STREAM[5],
               STREAM[4],STREAM[3],STREAM[2],STREAM[1],STREAM[0]}), .rd_data1 ({
               \$dummy [250],\$dummy [251],\$dummy [252],\$dummy [253],
               \$dummy [254],\$dummy [255],\$dummy [256],\$dummy [257]}), .addr1 (
               {FIFO_DEV_rtlc_wadd_n4[7],FIFO_DEV_rtlc_wadd_n4[6],
               FIFO_DEV_rtlc_wadd_n4[5],FIFO_DEV_rtlc_wadd_n4[4],
               FIFO_DEV_rtlc_wadd_n4[3],FIFO_DEV_rtlc_wadd_n4[2],
               FIFO_DEV_rtlc_wadd_n4[1],FIFO_DEV_rtlc_wadd_n4[0]}), .wr_clk1 (
               CLK_int), .rd_clk1 (\$dummy [258]), .wr_ena1 (\$dummy [259]), .rd_ena1 (
               \$dummy [260]), .ena1 (\$dummy [261]), .rst1 (\$dummy [262]), .regce1 (
               \$dummy [263]), .wr_data2 ({\$dummy [264],\$dummy [265],
               \$dummy [266],\$dummy [267],\$dummy [268],\$dummy [269],
               \$dummy [270],\$dummy [271]}), .rd_data2 ({nx12521z11,nx11524z4,
               nx10527z4,nx9530z4,nx8533z4,nx7536z4,nx6539z4,nx5542z4}), .addr2 (
               {FIFO_DEV_rtlc_radd_N1[7],FIFO_DEV_rtlc_radd_N1[6],
               FIFO_DEV_rtlc_radd_N1[5],FIFO_DEV_rtlc_radd_N1[4],
               FIFO_DEV_rtlc_radd_N1[3],FIFO_DEV_rtlc_radd_N1[2],
               FIFO_DEV_rtlc_radd_N1[1],FIFO_DEV_rtlc_radd_N1[0]}), .wr_clk2 (
               \$dummy [272]), .rd_clk2 (\$dummy [273]), .wr_ena2 (\$dummy [274]
               ), .rd_ena2 (\$dummy [275]), .ena2 (\$dummy [276]), .rst2 (
               \$dummy [277]), .regce2 (\$dummy [278]), .p_NOT_FIFO_DEV_rtlc5n43 (
               \$dummy [279]), .p_RST_int (RST_int), .p_NOT_CONDITION_0_ (
               NOT_CONDITION_0_), .p_WRITE (WRITE), .p_FIFO_DEV_rtlc_radd_N1_5___repl0 (
               FIFO_DEV_rtlc_radd_N1_5___repl0), .p_FIFO_DEV_rtlc_radd_N1_3___repl0 (
               FIFO_DEV_rtlc_radd_N1_3___repl0), .p_FIFO_DEV_rtlc_radd_N1_2___repl0 (
               FIFO_DEV_rtlc_radd_N1_2___repl0), .p_FIFO_DEV_rtlc_radd_N1_1___repl0 (
               FIFO_DEV_rtlc_radd_N1_1___repl0), .p_FIFO_DEV_rtlc_radd_N1_0___repl0 (
               FIFO_DEV_rtlc_radd_N1_0___repl0)) ;
    OUTBUF SIGN_REG_obuf_0_ (.PAD (SIGN_REG[0]), .D (SIGN_REG_dup_0[2])) ;
    OUTBUF SIGN_REG_obuf_1_ (.PAD (SIGN_REG[1]), .D (SIGN_REG_dup_0[3])) ;
    OUTBUF SIGN_REG_obuf_2_ (.PAD (SIGN_REG[2]), .D (SIGN_REG_dup_0[4])) ;
    OUTBUF SIGN_REG_obuf_3_ (.PAD (SIGN_REG[3]), .D (SIGN_REG_dup_0[5])) ;
    OUTBUF SIGN_REG_obuf_4_ (.PAD (SIGN_REG[4]), .D (SIGN_REG_dup_0[6])) ;
    OUTBUF SIGN_REG_obuf_5_ (.PAD (SIGN_REG[5]), .D (SIGN_REG_dup_0[7])) ;
    OUTBUF SIGN_REG_obuf_6_ (.PAD (SIGN_REG[6]), .D (SIGN_REG_dup_0[7])) ;
    OUTBUF SIGN_REG_obuf_7_ (.PAD (SIGN_REG[7]), .D (SIGN_REG_dup_0[7])) ;
    OUTBUF DATA_OUT_obuf_0_ (.PAD (DATA_OUT[0]), .D (DATA_OUT_dup_0[0])) ;
    OUTBUF DATA_OUT_obuf_1_ (.PAD (DATA_OUT[1]), .D (DATA_OUT_dup_0[1])) ;
    OUTBUF DATA_OUT_obuf_2_ (.PAD (DATA_OUT[2]), .D (DATA_OUT_dup_0[2])) ;
    OUTBUF DATA_OUT_obuf_3_ (.PAD (DATA_OUT[3]), .D (DATA_OUT_dup_0[3])) ;
    OUTBUF DATA_OUT_obuf_4_ (.PAD (DATA_OUT[4]), .D (DATA_OUT_dup_0[4])) ;
    OUTBUF DATA_OUT_obuf_5_ (.PAD (DATA_OUT[5]), .D (DATA_OUT_dup_0[5])) ;
    OUTBUF DATA_OUT_obuf_6_ (.PAD (DATA_OUT[6]), .D (DATA_OUT_dup_0[6])) ;
    OUTBUF DATA_OUT_obuf_7_ (.PAD (DATA_OUT[7]), .D (DATA_OUT_dup_0[7])) ;
    INBUF STB_KEY_ibuf (.Y (STB_KEY_int), .PAD (STB_KEY)) ;
    INBUF STB_DATA_ibuf (.Y (STB_DATA_int), .PAD (STB_DATA)) ;
    INBUF READ_ibuf (.Y (READ_int), .PAD (READ)) ;
    INBUF DATA_ibuf_0_ (.Y (DATA_int[0]), .PAD (DATA[0])) ;
    INBUF DATA_ibuf_1_ (.Y (DATA_int[1]), .PAD (DATA[1])) ;
    INBUF DATA_ibuf_2_ (.Y (DATA_int[2]), .PAD (DATA[2])) ;
    INBUF DATA_ibuf_3_ (.Y (DATA_int[3]), .PAD (DATA[3])) ;
    INBUF DATA_ibuf_4_ (.Y (DATA_int[4]), .PAD (DATA[4])) ;
    INBUF DATA_ibuf_5_ (.Y (DATA_int[5]), .PAD (DATA[5])) ;
    INBUF DATA_ibuf_6_ (.Y (DATA_int[6]), .PAD (DATA[6])) ;
    INBUF DATA_ibuf_7_ (.Y (DATA_int[7]), .PAD (DATA[7])) ;
    INBUF KEY_ibuf (.Y (KEY_int), .PAD (KEY)) ;
    DFN1 FIFO_DEV_ix12521z54533 (.Q (nx12521z6), .D (nx12521z3), .CLK (CLK_int)
         ) ;
    DFN1 FIFO_DEV_ix12521z54531 (.Q (nx12521z4), .D (nx12521z5), .CLK (CLK_int)
         ) ;
    DFN1 FIFO_DEV_ix11524z54529 (.Q (nx11524z2), .D (nx11524z1), .CLK (CLK_int)
         ) ;
    DFN1 FIFO_DEV_ix10527z54529 (.Q (nx10527z2), .D (nx10527z1), .CLK (CLK_int)
         ) ;
    DFN1 FIFO_DEV_ix9530z54529 (.Q (nx9530z2), .D (nx9530z1), .CLK (CLK_int)) ;
    DFN1 FIFO_DEV_ix8533z54529 (.Q (nx8533z2), .D (nx8533z1), .CLK (CLK_int)) ;
    DFN1 FIFO_DEV_ix7536z54529 (.Q (nx7536z2), .D (nx7536z1), .CLK (CLK_int)) ;
    DFN1 FIFO_DEV_ix6539z54529 (.Q (nx6539z2), .D (nx6539z1), .CLK (CLK_int)) ;
    DFN1 FIFO_DEV_ix5542z54529 (.Q (nx5542z2), .D (nx5542z1), .CLK (CLK_int)) ;
    DFN1 FIFO_DEV_ix12521z54535 (.Q (nx12521z8), .D (FIFO_DEV_not_dout_2n1s3), .CLK (
         CLK_int)) ;
    AND2 DATA_OUT_7__rename447 (.Y (DATA_OUT_dup_0[7]), .A (nx12521z1), .B (
         nx12521z3)) ;
    AND2 DATA_OUT_6__rename448 (.Y (DATA_OUT_dup_0[6]), .A (nx12521z1), .B (
         nx11524z1)) ;
    AND2 DATA_OUT_5__rename449 (.Y (DATA_OUT_dup_0[5]), .A (nx12521z1), .B (
         nx10527z1)) ;
    AND2 DATA_OUT_4__rename450 (.Y (DATA_OUT_dup_0[4]), .A (nx12521z1), .B (
         nx9530z1)) ;
    AND2 DATA_OUT_3__rename451 (.Y (DATA_OUT_dup_0[3]), .A (nx12521z1), .B (
         nx8533z1)) ;
    AND2 DATA_OUT_2__rename452 (.Y (DATA_OUT_dup_0[2]), .A (nx12521z1), .B (
         nx7536z1)) ;
    AND2 DATA_OUT_1__rename453 (.Y (DATA_OUT_dup_0[1]), .A (nx12521z1), .B (
         nx6539z1)) ;
    AND2 DATA_OUT_0__rename454 (.Y (DATA_OUT_dup_0[0]), .A (nx5542z1), .B (
         nx12521z1)) ;
    NAND3C CONDITION_1__rename455 (.Y (CONDITION_1_), .A (nx54297z1), .B (
           nx54297z3), .C (nx54297z4)) ;
    NAND3C NOT_CONDITION_0__rename456 (.Y (NOT_CONDITION_0_), .A (nx41852z1), .B (
           nx41852z3), .C (nx41852z4)) ;
    GND SIGN_REG_5__rename457 (.Y (SIGN_REG_dup_0[7])) ;
    XOR3 ENCR_DEV_t_1_0__rename458 (.Y (ENCR_DEV_t_1_0_), .A (nx13690z1), .B (
         ENCR_DEV_reg_str_1[65]), .C (ENCR_DEV_reg_str_1[92])) ;
    AX1C ENCR_DEV_t_1_1__rename459 (.Y (ENCR_DEV_t_1_1_), .A (
         ENCR_DEV_reg_str_1[90]), .B (ENCR_DEV_reg_str_1[89]), .C (nx12693z1)) ;
    AX1C ENCR_DEV_t_1_2__rename460 (.Y (ENCR_DEV_t_1_2_), .A (
         ENCR_DEV_reg_str_1[89]), .B (ENCR_DEV_reg_str_1[88]), .C (nx11696z1)) ;
    AX1C ENCR_DEV_t_1_3__rename461 (.Y (ENCR_DEV_t_1_3_), .A (
         ENCR_DEV_reg_str_1[88]), .B (ENCR_DEV_reg_str_1[87]), .C (nx10699z1)) ;
    AX1C ENCR_DEV_t_1_5__rename462 (.Y (ENCR_DEV_t_1_5_), .A (
         ENCR_DEV_reg_str_1[86]), .B (ENCR_DEV_reg_str_1[85]), .C (nx8705z1)) ;
    AX1C ENCR_DEV_t_1_6__rename463 (.Y (ENCR_DEV_t_1_6_), .A (
         ENCR_DEV_reg_str_1[85]), .B (ENCR_DEV_reg_str_1[84]), .C (nx7708z1)) ;
    XOR3 ENCR_DEV_t_2_0__rename464 (.Y (ENCR_DEV_t_2[0]), .A (nx22109z1), .B (
         ENCR_DEV_reg_str_2[68]), .C (ENCR_DEV_reg_str_2[83])) ;
    AX1C ENCR_DEV_t_2_1__rename465 (.Y (ENCR_DEV_t_2[1]), .A (
         ENCR_DEV_reg_str_2[81]), .B (ENCR_DEV_reg_str_2[80]), .C (nx21112z1)) ;
    AX1C ENCR_DEV_t_2_2__rename466 (.Y (ENCR_DEV_t_2[2]), .A (
         ENCR_DEV_reg_str_2[80]), .B (ENCR_DEV_reg_str_2[79]), .C (nx20115z1)) ;
    AX1C ENCR_DEV_t_2_3__rename467 (.Y (ENCR_DEV_t_2[3]), .A (
         ENCR_DEV_reg_str_2[79]), .B (ENCR_DEV_reg_str_2[78]), .C (nx19118z1)) ;
    AX1C ENCR_DEV_t_2_4__rename468 (.Y (ENCR_DEV_t_2[4]), .A (
         ENCR_DEV_reg_str_2[78]), .B (ENCR_DEV_reg_str_2[77]), .C (nx18121z1)) ;
    AX1C ENCR_DEV_t_2_5__rename469 (.Y (ENCR_DEV_t_2[5]), .A (
         ENCR_DEV_reg_str_2[77]), .B (ENCR_DEV_reg_str_2[76]), .C (nx17124z1)) ;
    AX1C ENCR_DEV_t_2_6__rename470 (.Y (ENCR_DEV_t_2[6]), .A (
         ENCR_DEV_reg_str_2[76]), .B (ENCR_DEV_reg_str_2[75]), .C (nx16127z1)) ;
    AX1C ENCR_DEV_t_2_7__rename471 (.Y (ENCR_DEV_t_2[7]), .A (
         ENCR_DEV_reg_str_2[75]), .B (ENCR_DEV_reg_str_2[74]), .C (nx15130z1)) ;
    XOR3 ENCR_DEV_t_3_0__rename472 (.Y (ENCR_DEV_t_3[0]), .A (nx35008z1), .B (
         ENCR_DEV_reg_str_3[65]), .C (ENCR_DEV_reg_str_3[110])) ;
    AX1C ENCR_DEV_t_3_1__rename473 (.Y (ENCR_DEV_t_3[1]), .A (
         ENCR_DEV_reg_str_3[108]), .B (ENCR_DEV_reg_str_3[107]), .C (nx36005z1)
         ) ;
    AX1C ENCR_DEV_t_3_2__rename474 (.Y (ENCR_DEV_t_3[2]), .A (
         ENCR_DEV_reg_str_3[107]), .B (ENCR_DEV_reg_str_3[106]), .C (nx37002z1)
         ) ;
    AX1C ENCR_DEV_t_3_3__rename475 (.Y (ENCR_DEV_t_3[3]), .A (
         ENCR_DEV_reg_str_3[106]), .B (ENCR_DEV_reg_str_3[105]), .C (nx37999z1)
         ) ;
    AX1C ENCR_DEV_t_3_4__rename476 (.Y (ENCR_DEV_t_3[4]), .A (
         ENCR_DEV_reg_str_3[105]), .B (ENCR_DEV_reg_str_3[104]), .C (nx38996z1)
         ) ;
    AX1C ENCR_DEV_t_3_5__rename477 (.Y (ENCR_DEV_t_3[5]), .A (
         ENCR_DEV_reg_str_3[104]), .B (ENCR_DEV_reg_str_3[103]), .C (nx39993z1)
         ) ;
    AX1C ENCR_DEV_t_3_6__rename478 (.Y (ENCR_DEV_t_3[6]), .A (
         ENCR_DEV_reg_str_3[103]), .B (ENCR_DEV_reg_str_3[102]), .C (nx40990z1)
         ) ;
    AX1C ENCR_DEV_t_3_7__rename479 (.Y (ENCR_DEV_t_3[7]), .A (
         ENCR_DEV_reg_str_3[102]), .B (ENCR_DEV_reg_str_3[101]), .C (nx41987z1)
         ) ;
    VCC ENCR_DEV_PWR_rename480 (.Y (ENCR_DEV_PWR)) ;
    NAND2B ENCR_DEV_ix7516z49935 (.Y (nx7516z2), .A (ENCR_DEV_prev[5]), .B (
           ENCR_DEV_prev_6__int)) ;
    NAND3C ENCR_DEV_ix3438z50934 (.Y (nx3438z3), .A (ENCR_DEV_prev[3]), .B (
           ENCR_DEV_prev[5]), .C (nx3438z4)) ;
    NAND2B ENCR_DEV_ix14495z49936 (.Y (nx14495z3), .A (ENCR_DEV_key_cnt[5]), .B (
           ENCR_DEV_key_cnt[4])) ;
    NAND3A NOT_ENCR_DEV_ix14495z50933 (.Y (nx14495z4), .A (nx43638z2), .B (
           ENCR_DEV_key_cnt[3]), .C (ENCR_DEV_key_cnt[2])) ;
    AO1C ENCR_DEV_ix14495z40558 (.Y (nx14495z2), .A (nx14495z3), .B (nx14495z4)
         , .C (ENCR_DEV_key_cnt[6])) ;
    NAND3C NOT_ENCR_DEV_ix15492z50936 (.Y (nx15492z5), .A (nx15492z6), .B (
           nx15492z7), .C (nx15492z8)) ;
    AO1C ENCR_DEV_ix15492z40559 (.Y (nx15492z3), .A (nx15492z4), .B (nx15492z5)
         , .C (ENCR_DEV_cnt_init[10])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_79__rename481 (.Y (
          ENCR_DEV_key_reg_12n5ss1[79]), .A (ENCR_DEV_prev[5]), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[78])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_78__rename482 (.Y (
          ENCR_DEV_key_reg_12n5ss1[78]), .A (ENCR_DEV_prev[5]), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[77])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_77__rename483 (.Y (
          ENCR_DEV_key_reg_12n5ss1[77]), .A (ENCR_DEV_prev[5]), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[76])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_76__rename484 (.Y (
          ENCR_DEV_key_reg_12n5ss1[76]), .A (ENCR_DEV_prev[5]), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[75])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_75__rename485 (.Y (
          ENCR_DEV_key_reg_12n5ss1[75]), .A (ENCR_DEV_prev[5]), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[74])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_74__rename486 (.Y (
          ENCR_DEV_key_reg_12n5ss1[74]), .A (ENCR_DEV_prev[5]), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[73])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_73__rename487 (.Y (
          ENCR_DEV_key_reg_12n5ss1[73]), .A (ENCR_DEV_prev[5]), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[72])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_72__rename488 (.Y (
          ENCR_DEV_key_reg_12n5ss1[72]), .A (ENCR_DEV_prev[5]), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[71])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_71__rename489 (.Y (
          ENCR_DEV_key_reg_12n5ss1[71]), .A (ENCR_DEV_prev[5]), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[70])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_70__rename490 (.Y (
          ENCR_DEV_key_reg_12n5ss1[70]), .A (ENCR_DEV_prev[5]), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[69])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_69__rename491 (.Y (
          ENCR_DEV_key_reg_12n5ss1[69]), .A (ENCR_DEV_prev[5]), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[68])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_68__rename492 (.Y (
          ENCR_DEV_key_reg_12n5ss1[68]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[67])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_67__rename493 (.Y (
          ENCR_DEV_key_reg_12n5ss1[67]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[66])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_66__rename494 (.Y (
          ENCR_DEV_key_reg_12n5ss1[66]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[65])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_65__rename495 (.Y (
          ENCR_DEV_key_reg_12n5ss1[65]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[64])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_64__rename496 (.Y (
          ENCR_DEV_key_reg_12n5ss1[64]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[63])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_63__rename497 (.Y (
          ENCR_DEV_key_reg_12n5ss1[63]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[62])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_62__rename498 (.Y (
          ENCR_DEV_key_reg_12n5ss1[62]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[61])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_61__rename499 (.Y (
          ENCR_DEV_key_reg_12n5ss1[61]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[60])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_60__rename500 (.Y (
          ENCR_DEV_key_reg_12n5ss1[60]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[59])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_59__rename501 (.Y (
          ENCR_DEV_key_reg_12n5ss1[59]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[58])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_58__rename502 (.Y (
          ENCR_DEV_key_reg_12n5ss1[58]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[57])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_57__rename503 (.Y (
          ENCR_DEV_key_reg_12n5ss1[57]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[56])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_56__rename504 (.Y (
          ENCR_DEV_key_reg_12n5ss1[56]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[55])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_55__rename505 (.Y (
          ENCR_DEV_key_reg_12n5ss1[55]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[54])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_54__rename506 (.Y (
          ENCR_DEV_key_reg_12n5ss1[54]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[53])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_53__rename507 (.Y (
          ENCR_DEV_key_reg_12n5ss1[53]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[52])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_52__rename508 (.Y (
          ENCR_DEV_key_reg_12n5ss1[52]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[51])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_51__rename509 (.Y (
          ENCR_DEV_key_reg_12n5ss1[51]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[50])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_50__rename510 (.Y (
          ENCR_DEV_key_reg_12n5ss1[50]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[49])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_49__rename511 (.Y (
          ENCR_DEV_key_reg_12n5ss1[49]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[48])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_48__rename512 (.Y (
          ENCR_DEV_key_reg_12n5ss1[48]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[47])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_47__rename513 (.Y (
          ENCR_DEV_key_reg_12n5ss1[47]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[46])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_46__rename514 (.Y (
          ENCR_DEV_key_reg_12n5ss1[46]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[45])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_45__rename515 (.Y (
          ENCR_DEV_key_reg_12n5ss1[45]), .A (ENCR_DEV_prev_5___repl2), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[44])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_44__rename516 (.Y (
          ENCR_DEV_key_reg_12n5ss1[44]), .A (ENCR_DEV_prev_5___repl1), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[43])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_43__rename517 (.Y (
          ENCR_DEV_key_reg_12n5ss1[43]), .A (ENCR_DEV_prev_5___repl1), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[42])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_42__rename518 (.Y (
          ENCR_DEV_key_reg_12n5ss1[42]), .A (ENCR_DEV_prev_5___repl1), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[41])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_41__rename519 (.Y (
          ENCR_DEV_key_reg_12n5ss1[41]), .A (ENCR_DEV_prev_5___repl1), .B (
          ENCR_DEV_prev_6__int), .C (ENCR_DEV_key_reg[40])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_40__rename520 (.Y (
          ENCR_DEV_key_reg_12n5ss1[40]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl1), .C (ENCR_DEV_key_reg[39])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_39__rename521 (.Y (
          ENCR_DEV_key_reg_12n5ss1[39]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl1), .C (ENCR_DEV_key_reg[38])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_38__rename522 (.Y (
          ENCR_DEV_key_reg_12n5ss1[38]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl1), .C (ENCR_DEV_key_reg[37])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_37__rename523 (.Y (
          ENCR_DEV_key_reg_12n5ss1[37]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl1), .C (ENCR_DEV_key_reg[36])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_36__rename524 (.Y (
          ENCR_DEV_key_reg_12n5ss1[36]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl1), .C (ENCR_DEV_key_reg[35])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_35__rename525 (.Y (
          ENCR_DEV_key_reg_12n5ss1[35]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl1), .C (ENCR_DEV_key_reg[34])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_34__rename526 (.Y (
          ENCR_DEV_key_reg_12n5ss1[34]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl1), .C (ENCR_DEV_key_reg[33])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_33__rename527 (.Y (
          ENCR_DEV_key_reg_12n5ss1[33]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl1), .C (ENCR_DEV_key_reg[32])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_32__rename528 (.Y (
          ENCR_DEV_key_reg_12n5ss1[32]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl1), .C (ENCR_DEV_key_reg[31])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_31__rename529 (.Y (
          ENCR_DEV_key_reg_12n5ss1[31]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl1), .C (ENCR_DEV_key_reg[30])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_30__rename530 (.Y (
          ENCR_DEV_key_reg_12n5ss1[30]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl1), .C (ENCR_DEV_key_reg[29])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_29__rename531 (.Y (
          ENCR_DEV_key_reg_12n5ss1[29]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl1), .C (ENCR_DEV_key_reg[28])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_28__rename532 (.Y (
          ENCR_DEV_key_reg_12n5ss1[28]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl1), .C (ENCR_DEV_key_reg[27])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_27__rename533 (.Y (
          ENCR_DEV_key_reg_12n5ss1[27]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl1), .C (ENCR_DEV_key_reg[26])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_26__rename534 (.Y (
          ENCR_DEV_key_reg_12n5ss1[26]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl1), .C (ENCR_DEV_key_reg[25])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_25__rename535 (.Y (
          ENCR_DEV_key_reg_12n5ss1[25]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl1), .C (ENCR_DEV_key_reg[24])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_24__rename536 (.Y (
          ENCR_DEV_key_reg_12n5ss1[24]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl1), .C (ENCR_DEV_key_reg[23])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_23__rename537 (.Y (
          ENCR_DEV_key_reg_12n5ss1[23]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl1), .C (ENCR_DEV_key_reg[22])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_22__rename538 (.Y (
          ENCR_DEV_key_reg_12n5ss1[22]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl1), .C (ENCR_DEV_key_reg[21])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_21__rename539 (.Y (
          ENCR_DEV_key_reg_12n5ss1[21]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl1), .C (ENCR_DEV_key_reg[20])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_20__rename540 (.Y (
          ENCR_DEV_key_reg_12n5ss1[20]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl0), .C (ENCR_DEV_key_reg[19])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_19__rename541 (.Y (
          ENCR_DEV_key_reg_12n5ss1[19]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl0), .C (ENCR_DEV_key_reg[18])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_18__rename542 (.Y (
          ENCR_DEV_key_reg_12n5ss1[18]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl0), .C (ENCR_DEV_key_reg[17])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_17__rename543 (.Y (
          ENCR_DEV_key_reg_12n5ss1[17]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl0), .C (ENCR_DEV_key_reg[16])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_16__rename544 (.Y (
          ENCR_DEV_key_reg_12n5ss1[16]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl0), .C (ENCR_DEV_key_reg[15])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_15__rename545 (.Y (
          ENCR_DEV_key_reg_12n5ss1[15]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl0), .C (ENCR_DEV_key_reg[14])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_14__rename546 (.Y (
          ENCR_DEV_key_reg_12n5ss1[14]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl0), .C (ENCR_DEV_key_reg[13])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_13__rename547 (.Y (
          ENCR_DEV_key_reg_12n5ss1[13]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl0), .C (ENCR_DEV_key_reg[12])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_12__rename548 (.Y (
          ENCR_DEV_key_reg_12n5ss1[12]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl0), .C (ENCR_DEV_key_reg[11])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_11__rename549 (.Y (
          ENCR_DEV_key_reg_12n5ss1[11]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl0), .C (ENCR_DEV_key_reg[10])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_10__rename550 (.Y (
          ENCR_DEV_key_reg_12n5ss1[10]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_5___repl0), .C (ENCR_DEV_key_reg[9])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_9__rename551 (.Y (ENCR_DEV_key_reg_12n5ss1[9]
          ), .A (ENCR_DEV_prev_6__int), .B (ENCR_DEV_prev_5___repl0), .C (
          ENCR_DEV_key_reg[8])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_8__rename552 (.Y (ENCR_DEV_key_reg_12n5ss1[8]
          ), .A (ENCR_DEV_prev_6__int), .B (ENCR_DEV_prev_5___repl0), .C (
          ENCR_DEV_key_reg[7])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_7__rename553 (.Y (ENCR_DEV_key_reg_12n5ss1[7]
          ), .A (ENCR_DEV_prev_6__int), .B (ENCR_DEV_prev_5___repl0), .C (
          ENCR_DEV_key_reg[6])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_6__rename554 (.Y (ENCR_DEV_key_reg_12n5ss1[6]
          ), .A (ENCR_DEV_prev_6__int), .B (ENCR_DEV_prev_5___repl0), .C (
          ENCR_DEV_key_reg[5])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_5__rename555 (.Y (ENCR_DEV_key_reg_12n5ss1[5]
          ), .A (ENCR_DEV_prev_6__int), .B (ENCR_DEV_prev_5___repl0), .C (
          ENCR_DEV_key_reg[4])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_4__rename556 (.Y (ENCR_DEV_key_reg_12n5ss1[4]
          ), .A (ENCR_DEV_prev_6__int), .B (ENCR_DEV_prev_5___repl0), .C (
          ENCR_DEV_key_reg[3])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_3__rename557 (.Y (ENCR_DEV_key_reg_12n5ss1[3]
          ), .A (ENCR_DEV_prev_6__int), .B (ENCR_DEV_prev_5___repl0), .C (
          ENCR_DEV_key_reg[2])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_2__rename558 (.Y (ENCR_DEV_key_reg_12n5ss1[2]
          ), .A (ENCR_DEV_prev_6__int), .B (ENCR_DEV_prev_5___repl0), .C (
          ENCR_DEV_key_reg[1])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_1__rename559 (.Y (ENCR_DEV_key_reg_12n5ss1[1]
          ), .A (ENCR_DEV_prev_6__int), .B (ENCR_DEV_prev_5___repl0), .C (
          ENCR_DEV_key_reg[0])) ;
    AND3B ENCR_DEV_key_reg_12n5ss1_0__rename560 (.Y (ENCR_DEV_key_reg_12n5ss1[0]
          ), .A (ENCR_DEV_prev_6__int), .B (ENCR_DEV_prev_5___repl0), .C (
          KEY_int)) ;
    NAND3C ENCR_DEV_rtlc12_X_0_n169_rename561 (.Y (ENCR_DEV_rtlc12_X_0_n169), .A (
           ENCR_DEV_prev_6__int), .B (ENCR_DEV_prev[7]), .C (
           ENCR_DEV_prev_5___repl0)) ;
    XA1 ENCR_DEV_stream_15n2ss1_7__rename562 (.Y (ENCR_DEV_stream_15n2ss1[7]), .A (
        nx41047z1), .B (nx41047z3), .C (nx1908z1)) ;
    XA1 ENCR_DEV_stream_15n2ss1_6__rename563 (.Y (ENCR_DEV_stream_15n2ss1[6]), .A (
        nx42044z1), .B (nx42044z3), .C (nx1908z1)) ;
    XA1 ENCR_DEV_stream_15n2ss1_5__rename564 (.Y (ENCR_DEV_stream_15n2ss1[5]), .A (
        nx43041z1), .B (nx43041z3), .C (nx1908z1)) ;
    XA1 ENCR_DEV_stream_15n2ss1_4__rename565 (.Y (ENCR_DEV_stream_15n2ss1[4]), .A (
        nx44038z1), .B (nx44038z3), .C (nx1908z1)) ;
    XA1 ENCR_DEV_stream_15n2ss1_3__rename566 (.Y (ENCR_DEV_stream_15n2ss1[3]), .A (
        nx45035z1), .B (nx45035z3), .C (nx1908z1)) ;
    XA1 ENCR_DEV_stream_15n2ss1_2__rename567 (.Y (ENCR_DEV_stream_15n2ss1[2]), .A (
        nx46032z1), .B (nx46032z3), .C (nx1908z1)) ;
    XA1 ENCR_DEV_stream_15n2ss1_1__rename568 (.Y (ENCR_DEV_stream_15n2ss1[1]), .A (
        nx47029z1), .B (nx47029z3), .C (nx1908z1)) ;
    XA1 ENCR_DEV_stream_15n2ss1_0__rename569 (.Y (ENCR_DEV_stream_15n2ss1[0]), .A (
        nx48026z1), .B (nx48026z3), .C (nx1908z1)) ;
    AND3B ENCR_DEV_reg_str_1_15n2ss1_92__rename570 (.Y (
          ENCR_DEV_reg_str_1_15n2ss1[92]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev[1]), .C (nx7977z1)) ;
    AND3B ENCR_DEV_reg_str_1_15n2ss1_91__rename571 (.Y (
          ENCR_DEV_reg_str_1_15n2ss1[91]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev[1]), .C (nx8974z1)) ;
    AND3B ENCR_DEV_reg_str_1_15n2ss1_90__rename572 (.Y (
          ENCR_DEV_reg_str_1_15n2ss1[90]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev[1]), .C (nx9971z1)) ;
    AND3B ENCR_DEV_reg_str_1_15n2ss1_89__rename573 (.Y (
          ENCR_DEV_reg_str_1_15n2ss1[89]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev[1]), .C (nx11967z1)) ;
    AND3B ENCR_DEV_reg_str_1_15n2ss1_88__rename574 (.Y (
          ENCR_DEV_reg_str_1_15n2ss1[88]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev[1]), .C (nx12964z1)) ;
    AND3B ENCR_DEV_reg_str_1_15n2ss1_87__rename575 (.Y (
          ENCR_DEV_reg_str_1_15n2ss1[87]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev[1]), .C (nx13961z1)) ;
    AND3B ENCR_DEV_reg_str_1_15n2ss1_86__rename576 (.Y (
          ENCR_DEV_reg_str_1_15n2ss1[86]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev[1]), .C (nx14958z1)) ;
    AND3B ENCR_DEV_reg_str_1_15n2ss1_85__rename577 (.Y (
          ENCR_DEV_reg_str_1_15n2ss1[85]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev[1]), .C (nx15955z1)) ;
    AND3B ENCR_DEV_reg_str_1_15n2ss1_84__rename578 (.Y (
          ENCR_DEV_reg_str_1_15n2ss1[84]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev[1]), .C (nx16952z1)) ;
    AND3B ENCR_DEV_reg_str_1_15n2ss1_83__rename579 (.Y (
          ENCR_DEV_reg_str_1_15n2ss1[83]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev[1]), .C (nx17949z1)) ;
    AND3B ENCR_DEV_reg_str_1_15n2ss1_82__rename580 (.Y (
          ENCR_DEV_reg_str_1_15n2ss1[82]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev[1]), .C (nx18946z1)) ;
    AND3B ENCR_DEV_reg_str_1_15n2ss1_81__rename581 (.Y (
          ENCR_DEV_reg_str_1_15n2ss1[81]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev[1]), .C (nx19943z1)) ;
    AND3B ENCR_DEV_reg_str_1_15n2ss1_80__rename582 (.Y (
          ENCR_DEV_reg_str_1_15n2ss1[80]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev[1]), .C (nx20940z1)) ;
    AND3B ENCR_DEV_reg_str_1_15n2ss1_79__rename583 (.Y (
          ENCR_DEV_reg_str_1_15n2ss1[79]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev[1]), .C (nx22936z1)) ;
    AND3B ENCR_DEV_reg_str_1_15n2ss1_78__rename584 (.Y (
          ENCR_DEV_reg_str_1_15n2ss1[78]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev[1]), .C (nx23933z1)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_77__rename585 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[77]), .A (nx24930z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx24930z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_76__rename586 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[76]), .A (nx25927z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx25927z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_75__rename587 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[75]), .A (nx26924z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx26924z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_74__rename588 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[74]), .A (nx27921z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx27921z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_73__rename589 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[73]), .A (nx28918z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx28918z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_72__rename590 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[72]), .A (nx29915z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx29915z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_71__rename591 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[71]), .A (nx30912z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx30912z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_70__rename592 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[70]), .A (nx31909z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx31909z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_69__rename593 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[69]), .A (nx33905z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx33905z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_68__rename594 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[68]), .A (nx34902z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx34902z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_67__rename595 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[67]), .A (nx35899z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx35899z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_66__rename596 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[66]), .A (nx36896z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx36896z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_65__rename597 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[65]), .A (nx37893z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx37893z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_64__rename598 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[64]), .A (nx38890z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx38890z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_63__rename599 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[63]), .A (nx39887z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx39887z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_62__rename600 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[62]), .A (nx40884z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx40884z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_61__rename601 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[61]), .A (nx41881z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx41881z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_60__rename602 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[60]), .A (nx42878z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx42878z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_59__rename603 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[59]), .A (nx44874z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx44874z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_58__rename604 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[58]), .A (nx45871z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx45871z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_57__rename605 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[57]), .A (nx46868z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx46868z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_56__rename606 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[56]), .A (nx47865z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx47865z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_55__rename607 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[55]), .A (nx48862z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx48862z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_54__rename608 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[54]), .A (nx49859z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx49859z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_53__rename609 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[53]), .A (nx50856z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx50856z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_52__rename610 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[52]), .A (nx51853z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx51853z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_51__rename611 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[51]), .A (nx52850z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx52850z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_50__rename612 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[50]), .A (nx53847z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx53847z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_49__rename613 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[49]), .A (nx55843z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx55843z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_48__rename614 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[48]), .A (nx56840z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx56840z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_47__rename615 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[47]), .A (nx57837z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx57837z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_46__rename616 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[46]), .A (nx58834z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx58834z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_45__rename617 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[45]), .A (nx59831z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx59831z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_44__rename618 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[44]), .A (nx60828z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx60828z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_43__rename619 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[43]), .A (nx61825z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx61825z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_42__rename620 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[42]), .A (nx62822z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx62822z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_41__rename621 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[41]), .A (nx63819z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx63819z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_40__rename622 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[40]), .A (nx64816z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx64816z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_39__rename623 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[39]), .A (nx1276z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx1276z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_38__rename624 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[38]), .A (nx2273z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx2273z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_37__rename625 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[37]), .A (nx3270z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx3270z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_36__rename626 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[36]), .A (nx4267z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx4267z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_35__rename627 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[35]), .A (nx5264z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx5264z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_34__rename628 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[34]), .A (nx6261z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx6261z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_33__rename629 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[33]), .A (nx7258z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx7258z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_32__rename630 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[32]), .A (nx8255z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx8255z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_31__rename631 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[31]), .A (nx9252z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx9252z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_30__rename632 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[30]), .A (nx10249z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx10249z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_29__rename633 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[29]), .A (nx12245z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx12245z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_28__rename634 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[28]), .A (nx13242z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx13242z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_27__rename635 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[27]), .A (nx14239z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx14239z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_26__rename636 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[26]), .A (nx15236z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx15236z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_25__rename637 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[25]), .A (nx16233z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx16233z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_24__rename638 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[24]), .A (nx17230z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx17230z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_23__rename639 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[23]), .A (nx18227z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx18227z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_22__rename640 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[22]), .A (nx19224z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx19224z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_21__rename641 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[21]), .A (nx20221z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx20221z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_20__rename642 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[20]), .A (nx21218z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx21218z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_19__rename643 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[19]), .A (nx23214z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx23214z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_18__rename644 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[18]), .A (nx24211z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx24211z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_17__rename645 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[17]), .A (nx25208z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx25208z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_16__rename646 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[16]), .A (nx26205z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx26205z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_15__rename647 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[15]), .A (nx27202z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx27202z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_14__rename648 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[14]), .A (nx28199z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx28199z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_13__rename649 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[13]), .A (nx29196z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx29196z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_12__rename650 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[12]), .A (nx30193z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx30193z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_11__rename651 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[11]), .A (nx31190z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx31190z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_10__rename652 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[10]), .A (nx32187z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx32187z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_9__rename653 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[9]), .A (nx44813z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx44813z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_8__rename654 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[8]), .A (nx43816z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx43816z2)) ;
    AO1C ENCR_DEV_reg_str_1_15n2ss1_7__rename655 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[7]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx42819z1), .C (nx42819z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_6__rename656 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[6]), .A (nx41822z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx41822z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_5__rename657 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[5]), .A (nx40825z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx40825z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_4__rename658 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[4]), .A (nx39828z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx39828z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_3__rename659 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[3]), .A (nx38831z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx38831z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_2__rename660 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[2]), .A (nx37834z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx37834z2)) ;
    MX2B ENCR_DEV_reg_str_1_15n2ss1_1__rename661 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[1]), .A (nx36837z1), .S (
         NOT_ENCR_DEV_rtlcn261_int), .B (nx36837z2)) ;
    AO1C ENCR_DEV_reg_str_1_15n2ss1_0__rename662 (.Y (
         ENCR_DEV_reg_str_1_15n2ss1[0]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx35840z1), .C (nx35840z2)) ;
    AND3B ENCR_DEV_reg_str_2_15n2ss1_83__rename663 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[83]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx61620z1)) ;
    AND3B ENCR_DEV_reg_str_2_15n2ss1_82__rename664 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[82]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx60623z1)) ;
    AND3B ENCR_DEV_reg_str_2_15n2ss1_81__rename665 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[81]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx59626z1)) ;
    AND3B ENCR_DEV_reg_str_2_15n2ss1_80__rename666 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[80]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx58629z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_79__rename667 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[79]), .A (nx56633z1), .B (
         NOT_ENCR_DEV_rtlcn261_int), .C (nx56633z2)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_78__rename668 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[78]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx55636z1), .C (nx55636z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_77__rename669 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[77]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx54639z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_76__rename670 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[76]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx53642z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_75__rename671 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[75]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx52645z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_74__rename672 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[74]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx51648z1), .C (nx51648z2)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_73__rename673 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[73]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx50651z1), .C (nx50651z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_72__rename674 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[72]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx49654z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_71__rename675 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[71]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx48657z1), .C (nx48657z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_70__rename676 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[70]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx47660z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_69__rename677 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[69]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx45664z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_68__rename678 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[68]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx44667z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_67__rename679 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[67]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx43670z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_66__rename680 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[66]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx42673z1), .C (nx42673z2)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_65__rename681 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[65]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx41676z1), .C (nx41676z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_64__rename682 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[64]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx40679z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_63__rename683 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[63]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx39682z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_62__rename684 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[62]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx38685z1), .C (nx38685z2)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_61__rename685 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[61]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx37688z2), .C (nx37688z3)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_60__rename686 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[60]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx36691z1), .C (nx36691z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_59__rename687 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[59]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx34695z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_58__rename688 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[58]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx33698z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_57__rename689 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[57]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx32701z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_56__rename690 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[56]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx31704z1), .C (nx31704z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_55__rename691 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[55]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx30707z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_54__rename692 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[54]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx29710z1), .C (nx29710z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_53__rename693 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[53]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx28713z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_52__rename694 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[52]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx27716z1), .C (nx27716z2)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_51__rename695 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[51]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx26719z1), .C (nx26719z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_50__rename696 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[50]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx25722z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_49__rename697 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[49]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx23726z1), .C (nx23726z2)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_48__rename698 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[48]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx22729z1), .C (nx22729z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_47__rename699 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[47]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx21732z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_46__rename700 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[46]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx20735z1), .C (nx20735z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_45__rename701 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[45]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx19738z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_44__rename702 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[44]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx18741z1), .C (nx18741z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_43__rename703 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[43]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx17744z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_42__rename704 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[42]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx16747z1), .C (nx16747z2)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_41__rename705 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[41]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx15750z1), .C (nx15750z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_40__rename706 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[40]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx14753z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_39__rename707 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[39]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx12757z1), .C (nx12757z2)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_38__rename708 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[38]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx11760z1), .C (nx11760z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_37__rename709 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[37]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx10763z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_36__rename710 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[36]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx9766z1), .C (nx9766z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_35__rename711 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[35]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx8769z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_34__rename712 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[34]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx7772z1), .C (nx7772z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_33__rename713 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[33]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx6775z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_32__rename714 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[32]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx5778z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_31__rename715 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[31]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx4781z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_30__rename716 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[30]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx3784z1), .C (nx3784z2)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_29__rename717 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[29]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx1788z1), .C (nx1788z2)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_28__rename718 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[28]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx791z1), .C (nx791z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_27__rename719 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[27]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx65330z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_26__rename720 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[26]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx64333z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_25__rename721 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[25]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx63336z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_24__rename722 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[24]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx62339z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_23__rename723 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[23]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx61342z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_22__rename724 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[22]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx60345z1), .C (nx60345z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_21__rename725 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[21]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx59348z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_20__rename726 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[20]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx58351z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_19__rename727 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[19]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx56355z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_18__rename728 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[18]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx55358z1), .C (nx55358z2)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_17__rename729 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[17]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx54361z1), .C (nx54361z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_16__rename730 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[16]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx53364z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_15__rename731 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[15]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx52367z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_14__rename732 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[14]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx51370z1), .C (nx51370z2)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_13__rename733 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[13]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx50373z1), .C (nx50373z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_12__rename734 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[12]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx49376z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_11__rename735 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[11]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx48379z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_10__rename736 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[10]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx47382z1), .C (nx47382z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_9__rename737 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[9]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx16502z1)) ;
    AO1E ENCR_DEV_reg_str_2_15n2ss1_8__rename738 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[8]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx17499z1), .C (nx17499z2)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_7__rename739 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[7]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx18496z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_6__rename740 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[6]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx19493z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_5__rename741 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[5]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx20490z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_4__rename742 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[4]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx21487z1)) ;
    AO1C ENCR_DEV_reg_str_2_15n2ss1_3__rename743 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[3]), .A (b_0__int), .B (nx22484z1), .C (
         nx22484z3)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_2__rename744 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[2]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx23481z1)) ;
    AND2A ENCR_DEV_reg_str_2_15n2ss1_1__rename745 (.Y (
          ENCR_DEV_reg_str_2_15n2ss1[1]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
          nx24478z1)) ;
    AO1C ENCR_DEV_reg_str_2_15n2ss1_0__rename746 (.Y (
         ENCR_DEV_reg_str_2_15n2ss1[0]), .A (b_0__int), .B (nx25475z1), .C (
         nx25475z3)) ;
    AO1E ENCR_DEV_reg_str_3_15n2ss1_110__rename747 (.Y (
         ENCR_DEV_reg_str_3_15n2ss1[110]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx38120z1), .C (nx38120z2)) ;
    AO1E ENCR_DEV_reg_str_3_15n2ss1_109__rename748 (.Y (
         ENCR_DEV_reg_str_3_15n2ss1[109]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx36124z1), .C (nx36124z2)) ;
    AO1E ENCR_DEV_reg_str_3_15n2ss1_108__rename749 (.Y (
         ENCR_DEV_reg_str_3_15n2ss1[108]), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         nx35127z1), .C (nx35127z2)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_107__rename750 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[107]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx34130z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_106__rename751 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[106]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx33133z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_105__rename752 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[105]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx32136z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_104__rename753 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[104]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx31139z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_103__rename754 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[103]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx30142z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_102__rename755 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[102]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx29145z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_101__rename756 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[101]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx28148z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_100__rename757 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[100]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx27151z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_99__rename758 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[99]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx38468z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_98__rename759 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[98]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx39465z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_97__rename760 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[97]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx40462z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_96__rename761 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[96]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx41459z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_95__rename762 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[95]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx42456z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_94__rename763 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[94]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx43453z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_93__rename764 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[93]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx44450z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_92__rename765 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[92]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx45447z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_91__rename766 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[91]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx46444z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_90__rename767 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[90]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx47441z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_89__rename768 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[89]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx49437z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_88__rename769 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[88]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl4), .C (nx50434z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_87__rename770 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[87]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx51431z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_86__rename771 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[86]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx52428z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_85__rename772 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[85]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx53425z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_84__rename773 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[84]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx54422z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_83__rename774 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[83]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx55419z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_82__rename775 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[82]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx56416z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_81__rename776 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[81]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx57413z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_80__rename777 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[80]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx58410z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_79__rename778 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[79]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx60406z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_78__rename779 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[78]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx61403z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_77__rename780 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[77]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx62400z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_76__rename781 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[76]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx63397z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_75__rename782 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[75]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx64394z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_74__rename783 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[74]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx65391z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_73__rename784 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[73]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx852z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_72__rename785 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[72]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx1849z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_71__rename786 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[71]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx2846z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_70__rename787 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[70]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx3843z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_69__rename788 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[69]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx5839z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_68__rename789 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[68]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx6836z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_67__rename790 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[67]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx7833z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_66__rename791 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[66]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx8830z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_65__rename792 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[65]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx9827z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_64__rename793 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[64]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl3), .C (nx10824z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_63__rename794 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[63]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx11821z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_62__rename795 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[62]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx12818z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_61__rename796 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[61]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx13815z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_60__rename797 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[60]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx14812z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_59__rename798 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[59]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx16808z2)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_58__rename799 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[58]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx17805z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_57__rename800 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[57]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx18802z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_56__rename801 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[56]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx19799z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_55__rename802 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[55]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx20796z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_54__rename803 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[54]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx21793z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_53__rename804 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[53]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx22790z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_52__rename805 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[52]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx23787z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_51__rename806 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[51]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx24784z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_50__rename807 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[50]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx25781z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_49__rename808 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[49]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx27777z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_48__rename809 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[48]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx28774z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_47__rename810 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[47]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx29771z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_46__rename811 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[46]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx30768z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_45__rename812 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[45]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx31765z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_44__rename813 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[44]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx32762z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_43__rename814 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[43]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx33759z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_42__rename815 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[42]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx34756z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_41__rename816 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[41]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx35753z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_40__rename817 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[40]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl2), .C (nx36750z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_39__rename818 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[39]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx38746z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_38__rename819 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[38]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx39743z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_37__rename820 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[37]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx40740z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_36__rename821 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[36]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx41737z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_35__rename822 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[35]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx42734z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_34__rename823 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[34]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx43731z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_33__rename824 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[33]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx44728z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_32__rename825 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[32]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx45725z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_31__rename826 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[31]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx46722z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_30__rename827 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[30]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx47719z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_29__rename828 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[29]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx49715z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_28__rename829 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[28]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx50712z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_27__rename830 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[27]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx51709z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_26__rename831 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[26]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx52706z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_25__rename832 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[25]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx53703z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_24__rename833 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[24]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx54700z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_23__rename834 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[23]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx55697z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_22__rename835 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[22]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx56694z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_21__rename836 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[21]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx57691z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_20__rename837 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[20]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx58688z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_19__rename838 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[19]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx60684z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_18__rename839 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[18]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx61681z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_17__rename840 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[17]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx62678z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_16__rename841 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[16]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl1), .C (nx63675z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_15__rename842 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[15]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl0), .C (nx64672z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_14__rename843 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[14]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl0), .C (nx133z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_13__rename844 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[13]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl0), .C (nx1130z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_12__rename845 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[12]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl0), .C (nx2127z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_11__rename846 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[11]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl0), .C (nx3124z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_10__rename847 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[10]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl0), .C (nx4121z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_9__rename848 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[9]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl0), .C (nx12281z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_8__rename849 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[8]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl0), .C (nx13278z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_7__rename850 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[7]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl0), .C (nx14275z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_6__rename851 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[6]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl0), .C (nx15272z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_5__rename852 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[5]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl0), .C (nx16269z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_4__rename853 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[4]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl0), .C (nx17266z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_3__rename854 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[3]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl0), .C (nx18263z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_2__rename855 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[2]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl0), .C (nx19260z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_1__rename856 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[1]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl0), .C (nx20257z1)) ;
    AND3B ENCR_DEV_reg_str_3_15n2ss1_0__rename857 (.Y (
          ENCR_DEV_reg_str_3_15n2ss1[0]), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev_1___repl0), .C (nx21254z1)) ;
    NAND2B ENCR_DEV_ix8587z49934 (.Y (nx8587z1), .A (ENCR_DEV_prev_6__int), .B (
           ENCR_DEV_prev[2])) ;
    NAND2B ENCR_DEV_ix63528z49934 (.Y (nx63528z1), .A (ENCR_DEV_prev_6__int), .B (
           ENCR_DEV_prev[3])) ;
    AND3C ENCR_DEV_ix46110z2958 (.Y (nx46110z1), .A (ENCR_DEV_prev_6__int), .B (
          ENCR_DEV_prev[2]), .C (ENCR_DEV_prev[3])) ;
    NAND2 NOT_ENCR_DEV_t_1_4_16n1s20_rename858 (.Y (NOT_ENCR_DEV_t_1_4_16n1s20)
          , .A (ENCR_DEV_reg_str_1[87]), .B (ENCR_DEV_reg_str_1[86])) ;
    NAND2 NOT_ENCR_DEV_t_1_7_16n1s32_rename859 (.Y (NOT_ENCR_DEV_t_1_7_16n1s32)
          , .A (ENCR_DEV_reg_str_1[84]), .B (ENCR_DEV_reg_str_1[83])) ;
    NAND3C ENCR_DEV_ix18636z50932 (.Y (nx18636z1), .A (ENCR_DEV_prev[7]), .B (
           ENCR_DEV_prev[4]), .C (ENCR_DEV_prev[2])) ;
    AND2 ENCR_DEV_ix1908z48514 (.Y (nx1908z1), .A (ENCR_DEV_strob_data_tmp), .B (
         ENCR_DEV_prev[2])) ;
    AO1C ENCR_DEV_ix10507z40557 (.Y (nx10507z1), .A (nx10507z2), .B (nx10507z3)
         , .C (nx10507z5)) ;
    AO1A ENCR_DEV_ix9510z40555 (.Y (nx9510z1), .A (nx9510z2), .B (nx10507z3), .C (
         nx9510z8)) ;
    AOI1A ENCR_DEV_ix15492z47388 (.Y (nx15492z1), .A (ENCR_DEV_prev[7]), .B (
          nx15492z2), .C (STB_KEY_int)) ;
    AO1C ENCR_DEV_ix36622z40557 (.Y (nx36622z1), .A (nx36622z2), .B (nx14495z2)
         , .C (nx36622z3)) ;
    AND2 ENCR_DEV_ix13498z48514 (.Y (nx13498z1), .A (ENCR_DEV_prev[4]), .B (
         STB_DATA_int)) ;
    AO1E ENCR_DEV_ix11504z40559 (.Y (nx11504z1), .A (nx11504z2), .B (nx11504z18)
         , .C (nx11504z22)) ;
    AO1A ENCR_DEV_ix7516z40555 (.Y (nx7516z1), .A (STB_KEY_int), .B (
         ENCR_DEV_prev[0]), .C (nx7516z2)) ;
    AND3B ENCR_DEV_ix3438z2957 (.Y (nx3438z1), .A (nx3438z2), .B (nx3438z3), .C (
          nx3438z5)) ;
    NAND2A ENCR_DEV_ix3438z49937 (.Y (nx3438z5), .A (nx14495z2), .B (
           ENCR_DEV_prev_1___repl0)) ;
    NAND2 NOT_ENCR_DEV_ix10507z24342 (.Y (nx10507z5), .A (CONDITION_1_), .B (
          ENCR_DEV_prev[3])) ;
    AO1A NOT_ENCR_DEV_ix9510z40563 (.Y (nx9510z9), .A (ENCR_DEV_cnt_init[11]), .B (
         nx15492z3), .C (nx9510z10)) ;
    NAND3A NOT_ENCR_DEV_ix15492z50931 (.Y (nx15492z2), .A (ENCR_DEV_cnt_init[11]
           ), .B (nx15492z3), .C (ENCR_DEV_prev[8])) ;
    AO1C NOT_ENCR_DEV_ix36622z40559 (.Y (nx36622z3), .A (ENCR_DEV_prev[8]), .B (
         nx3438z5), .C (STB_KEY_int)) ;
    NAND3B NOT_ENCR_DEV_ix11504z50953 (.Y (nx11504z22), .A (STB_KEY_int), .B (
           STB_DATA_int), .C (ENCR_DEV_prev[4])) ;
    NAND3 ENCR_DEV_ix45632z24339 (.Y (nx45632z3), .A (nx14495z3), .B (
          ENCR_DEV_key_cnt[6]), .C (ENCR_DEV_prev_1___repl0)) ;
    AND2A ENCR_DEV_ix25368z1959 (.Y (nx25368z1), .A (ENCR_DEV_strob_data_tmp), .B (
          ENCR_DEV_prev[2])) ;
    NAND3B NOT_ENCR_DEV_ix9510z50933 (.Y (nx9510z3), .A (nx9510z4), .B (nx9510z6
           ), .C (ENCR_DEV_encry_cnt[0])) ;
    NAND3C NOT_ENCR_DEV_ix10507z50934 (.Y (nx10507z3), .A (nx10507z4), .B (
           nx11504z10), .C (nx11504z19)) ;
    AX1C ENCR_DEV_ix35008z8206 (.Y (nx35008z1), .A (ENCR_DEV_reg_str_3[109]), .B (
         ENCR_DEV_reg_str_3[108]), .C (ENCR_DEV_reg_str_1[68])) ;
    AX1C ENCR_DEV_ix13690z8206 (.Y (nx13690z1), .A (ENCR_DEV_reg_str_1[91]), .B (
         ENCR_DEV_reg_str_1[90]), .C (ENCR_DEV_reg_str_2[77])) ;
    XOR3 ENCR_DEV_ix16127z10877 (.Y (nx16127z1), .A (ENCR_DEV_reg_str_2[77]), .B (
         ENCR_DEV_reg_str_2[62]), .C (ENCR_DEV_reg_str_3[80])) ;
    XOR3 ENCR_DEV_ix37999z10877 (.Y (nx37999z1), .A (ENCR_DEV_reg_str_3[107]), .B (
         ENCR_DEV_reg_str_1[65]), .C (ENCR_DEV_reg_str_3[62])) ;
    AX1C ENCR_DEV_ix22109z8206 (.Y (nx22109z1), .A (ENCR_DEV_reg_str_2[82]), .B (
         ENCR_DEV_reg_str_2[81]), .C (ENCR_DEV_reg_str_3[86])) ;
    XOR3 ENCR_DEV_ix36005z10877 (.Y (nx36005z1), .A (ENCR_DEV_reg_str_3[109]), .B (
         ENCR_DEV_reg_str_3[64]), .C (ENCR_DEV_reg_str_1[67])) ;
    XOR3 ENCR_DEV_ix21112z10877 (.Y (nx21112z1), .A (ENCR_DEV_reg_str_2[82]), .B (
         ENCR_DEV_reg_str_2[67]), .C (ENCR_DEV_reg_str_3[85])) ;
    XOR3 ENCR_DEV_ix12693z10877 (.Y (nx12693z1), .A (ENCR_DEV_reg_str_1[91]), .B (
         ENCR_DEV_reg_str_1[64]), .C (ENCR_DEV_reg_str_2[76])) ;
    XOR3 ENCR_DEV_ix38996z10877 (.Y (nx38996z1), .A (ENCR_DEV_reg_str_3[106]), .B (
         ENCR_DEV_reg_str_1[64]), .C (ENCR_DEV_reg_str_3[61])) ;
    XOR3 ENCR_DEV_ix37002z10877 (.Y (nx37002z1), .A (ENCR_DEV_reg_str_3[108]), .B (
         ENCR_DEV_reg_str_3[63]), .C (ENCR_DEV_reg_str_1[66])) ;
    XOR3 ENCR_DEV_ix20115z10877 (.Y (nx20115z1), .A (ENCR_DEV_reg_str_2[81]), .B (
         ENCR_DEV_reg_str_2[66]), .C (ENCR_DEV_reg_str_3[84])) ;
    XOR3 ENCR_DEV_ix11696z10877 (.Y (nx11696z1), .A (ENCR_DEV_reg_str_1[90]), .B (
         ENCR_DEV_reg_str_1[63]), .C (ENCR_DEV_reg_str_2[75])) ;
    XOR3 ENCR_DEV_ix39993z10877 (.Y (nx39993z1), .A (ENCR_DEV_reg_str_3[105]), .B (
         ENCR_DEV_reg_str_1[63]), .C (ENCR_DEV_reg_str_3[60])) ;
    XOR3 ENCR_DEV_ix19118z10877 (.Y (nx19118z1), .A (ENCR_DEV_reg_str_2[80]), .B (
         ENCR_DEV_reg_str_2[65]), .C (ENCR_DEV_reg_str_3[83])) ;
    XOR3 ENCR_DEV_ix10699z10877 (.Y (nx10699z1), .A (ENCR_DEV_reg_str_1[89]), .B (
         ENCR_DEV_reg_str_1[62]), .C (ENCR_DEV_reg_str_2[74])) ;
    XOR3 ENCR_DEV_ix40990z10877 (.Y (nx40990z1), .A (ENCR_DEV_reg_str_3[104]), .B (
         ENCR_DEV_reg_str_1[62]), .C (ENCR_DEV_reg_str_3[59])) ;
    XOR3 ENCR_DEV_ix18121z10877 (.Y (nx18121z1), .A (ENCR_DEV_reg_str_2[79]), .B (
         ENCR_DEV_reg_str_2[64]), .C (ENCR_DEV_reg_str_3[82])) ;
    XOR3 ENCR_DEV_ix22484z10878 (.Y (nx22484z2), .A (ENCR_DEV_reg_str_1[88]), .B (
         ENCR_DEV_reg_str_1[61]), .C (ENCR_DEV_reg_str_2[73])) ;
    XOR3 ENCR_DEV_ix41987z10877 (.Y (nx41987z1), .A (ENCR_DEV_reg_str_3[103]), .B (
         ENCR_DEV_reg_str_1[61]), .C (ENCR_DEV_reg_str_3[58])) ;
    XOR3 ENCR_DEV_ix17124z10877 (.Y (nx17124z1), .A (ENCR_DEV_reg_str_2[78]), .B (
         ENCR_DEV_reg_str_2[63]), .C (ENCR_DEV_reg_str_3[81])) ;
    XOR3 ENCR_DEV_ix8705z10877 (.Y (nx8705z1), .A (ENCR_DEV_reg_str_1[87]), .B (
         ENCR_DEV_reg_str_1[60]), .C (ENCR_DEV_reg_str_2[72])) ;
    XOR3 ENCR_DEV_ix7708z10877 (.Y (nx7708z1), .A (ENCR_DEV_reg_str_1[86]), .B (
         ENCR_DEV_reg_str_1[59]), .C (ENCR_DEV_reg_str_2[71])) ;
    XOR3 ENCR_DEV_ix15130z10877 (.Y (nx15130z1), .A (ENCR_DEV_reg_str_2[76]), .B (
         ENCR_DEV_reg_str_2[61]), .C (ENCR_DEV_reg_str_3[79])) ;
    XOR3 ENCR_DEV_ix25475z10878 (.Y (nx25475z2), .A (ENCR_DEV_reg_str_1[85]), .B (
         ENCR_DEV_reg_str_1[58]), .C (ENCR_DEV_reg_str_2[70])) ;
    NAND2 NOT_FIFO_DEV_ix32158z24340 (.Y (nx32158z2), .A (NOT_CONDITION_0_), .B (
          WRITE)) ;
    INV FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_0__rename860 (.Y (
        FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_0_), .A (
        FIFO_DEV_rtlc_radd_N1_0___repl0)) ;
    AX1C FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_2__rename861 (.Y (
         FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_2_), .A (
         FIFO_DEV_rtlc_radd_N1_1___repl0), .B (FIFO_DEV_rtlc_radd_N1_0___repl0)
         , .C (FIFO_DEV_rtlc_radd_N1_2___repl0)) ;
    AX1 FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_3__rename862 (.Y (
        FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_3_), .A (nx4093z3), .B (
        FIFO_DEV_rtlc_radd_N1_2___repl0), .C (FIFO_DEV_rtlc_radd_N1_3___repl0)
        ) ;
    XNOR2 FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_4__rename863 (.Y (
          FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_4_), .A (nx4093z2), .B (
          FIFO_DEV_rtlc_radd_N1[4])) ;
    AX1 FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_5__rename864 (.Y (
        FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_5_), .A (nx4093z2), .B (
        FIFO_DEV_rtlc_radd_N1[4]), .C (FIFO_DEV_rtlc_radd_N1_5___repl0)) ;
    XNOR2 FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_6__rename865 (.Y (
          FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_6_), .A (nx4093z1), .B (
          FIFO_DEV_rtlc_radd_N1[6])) ;
    AX1 FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_7__rename866 (.Y (
        FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_7_), .A (nx4093z1), .B (
        FIFO_DEV_rtlc_radd_N1[6]), .C (FIFO_DEV_rtlc_radd_N1[7])) ;
    NAND2 NOT_FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_ix4093z24340 (.Y (
          nx4093z3), .A (FIFO_DEV_rtlc_radd_N1_1___repl0), .B (
          FIFO_DEV_rtlc_radd_N1_0___repl0)) ;
    NAND3A NOT_FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_ix4093z50931 (.Y (
           nx4093z2), .A (nx4093z3), .B (FIFO_DEV_rtlc_radd_N1_2___repl0), .C (
           FIFO_DEV_rtlc_radd_N1_3___repl0)) ;
    NAND3A NOT_FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_ix4093z50930 (.Y (
           nx4093z1), .A (nx4093z2), .B (FIFO_DEV_rtlc_radd_N1[4]), .C (
           FIFO_DEV_rtlc_radd_N1_5___repl0)) ;
    AO1C FIFO_DEV_ix12521z40559 (.Y (nx12521z3), .A (nx12521z4), .B (nx12521z6)
         , .C (nx12521z7)) ;
    AO1C FIFO_DEV_ix11524z40557 (.Y (nx11524z1), .A (nx12521z4), .B (nx11524z2)
         , .C (nx11524z3)) ;
    AO1C FIFO_DEV_ix10527z40557 (.Y (nx10527z1), .A (nx12521z4), .B (nx10527z2)
         , .C (nx10527z3)) ;
    AO1C FIFO_DEV_ix9530z40557 (.Y (nx9530z1), .A (nx12521z4), .B (nx9530z2), .C (
         nx9530z3)) ;
    AO1C FIFO_DEV_ix8533z40557 (.Y (nx8533z1), .A (nx12521z4), .B (nx8533z2), .C (
         nx8533z3)) ;
    AO1C FIFO_DEV_ix7536z40557 (.Y (nx7536z1), .A (nx12521z4), .B (nx7536z2), .C (
         nx7536z3)) ;
    AO1C FIFO_DEV_ix6539z40557 (.Y (nx6539z1), .A (nx12521z4), .B (nx6539z2), .C (
         nx6539z3)) ;
    AO1C FIFO_DEV_ix5542z40557 (.Y (nx5542z1), .A (nx12521z4), .B (nx5542z2), .C (
         nx5542z3)) ;
    NAND3C b_0__rename867 (.Y (b_0_), .A (ENCR_DEV_prev_6__int), .B (
           ENCR_DEV_prev_1___repl0), .C (ENCR_DEV_prev_8___repl0)) ;
    NAND3C NOT_ENCR_DEV_ix37688z50933 (.Y (nx37688z1), .A (ENCR_DEV_prev_6__int)
           , .B (ENCR_DEV_prev_1___repl0), .C (ENCR_DEV_prev[7])) ;
    XA1B sclear_and_0_dup_147_rename868 (.Y (sclear_and_0_dup_147), .A (
         ENCR_DEV_cnt_init[0]), .B (ENCR_DEV_prev[8]), .C (nx8587z1)) ;
    XA1C sclear_and_1_dup_148_rename869 (.Y (sclear_and_1_dup_148), .A (
         nx27756z1), .B (ENCR_DEV_cnt_init[1]), .C (nx8587z1)) ;
    XA1C sclear_and_2_dup_149_rename870 (.Y (sclear_and_2_dup_149), .A (
         nx61539z3), .B (ENCR_DEV_cnt_init[2]), .C (nx8587z1)) ;
    AND3B sclear_and_3_dup_150_rename871 (.Y (sclear_and_3_dup_150), .A (
          ENCR_DEV_prev_6__int), .B (ENCR_DEV_prev[2]), .C (inc_d_3_)) ;
    XA1C sclear_and_4_dup_151_rename872 (.Y (sclear_and_4_dup_151), .A (
         nx61539z2), .B (ENCR_DEV_cnt_init[4]), .C (nx8587z1)) ;
    AND3B sclear_and_5_dup_152_rename873 (.Y (sclear_and_5_dup_152), .A (
          ENCR_DEV_prev_6__int), .B (ENCR_DEV_prev[2]), .C (inc_d_5_)) ;
    XA1C sclear_and_6_dup_153_rename874 (.Y (sclear_and_6_dup_153), .A (
         ENCR_DEV_cnt_init[6]), .B (nx54095z1), .C (nx8587z1)) ;
    XA1C sclear_and_7_dup_154_rename875 (.Y (sclear_and_7_dup_154), .A (
         ENCR_DEV_cnt_init[7]), .B (nx34195z1), .C (nx8587z1)) ;
    XA1C sclear_and_8_dup_155_rename876 (.Y (sclear_and_8_dup_155), .A (
         ENCR_DEV_cnt_init[8]), .B (nx61539z1), .C (nx8587z1)) ;
    AND3B sclear_and_9_dup_156_rename877 (.Y (sclear_and_9_dup_156), .A (
          ENCR_DEV_prev_6__int), .B (ENCR_DEV_prev[2]), .C (inc_d_9_)) ;
    XA1C sclear_and_10_dup_157_rename878 (.Y (sclear_and_10_dup_157), .A (
         ENCR_DEV_cnt_init[10]), .B (nx8464z1), .C (nx8587z1)) ;
    XA1C sclear_and_11_dup_158_rename879 (.Y (sclear_and_11_dup_158), .A (
         nx34318z1), .B (ENCR_DEV_cnt_init[11]), .C (nx8587z1)) ;
    NAND2 NOT_ix34195z24339 (.Y (nx34195z2), .A (ENCR_DEV_cnt_init[5]), .B (
          ENCR_DEV_cnt_init[4])) ;
    NAND2 NOT_ix34318z24339 (.Y (nx34318z2), .A (ENCR_DEV_cnt_init[9]), .B (
          ENCR_DEV_cnt_init[8])) ;
    NAND2 NOT_ix27756z24338 (.Y (nx27756z1), .A (ENCR_DEV_cnt_init[0]), .B (
          ENCR_DEV_prev[8])) ;
    NAND3 NOT_ix61539z24339 (.Y (nx61539z3), .A (ENCR_DEV_cnt_init[0]), .B (
          ENCR_DEV_prev[8]), .C (ENCR_DEV_cnt_init[1])) ;
    NAND2 NOT_ix61539z24341 (.Y (nx61539z4), .A (ENCR_DEV_cnt_init[7]), .B (
          ENCR_DEV_cnt_init[6])) ;
    NAND3A NOT_ix61539z50931 (.Y (nx61539z2), .A (nx61539z3), .B (
           ENCR_DEV_cnt_init[3]), .C (ENCR_DEV_cnt_init[2])) ;
    NAND3A NOT_ix54095z50930 (.Y (nx54095z1), .A (nx61539z2), .B (
           ENCR_DEV_cnt_init[5]), .C (ENCR_DEV_cnt_init[4])) ;
    NAND3C NOT_ix61539z50932 (.Y (nx61539z1), .A (nx61539z2), .B (nx34195z2), .C (
           nx61539z4)) ;
    NAND3B NOT_ix34195z50931 (.Y (nx34195z1), .A (nx61539z2), .B (nx34195z2), .C (
           ENCR_DEV_cnt_init[6])) ;
    NAND3A NOT_ix8464z50930 (.Y (nx8464z1), .A (nx61539z1), .B (
           ENCR_DEV_cnt_init[9]), .C (ENCR_DEV_cnt_init[8])) ;
    NAND3B NOT_ix34318z50931 (.Y (nx34318z1), .A (nx34318z2), .B (nx61539z1), .C (
           ENCR_DEV_cnt_init[10])) ;
    AX1 inc_d_3__rename880 (.Y (inc_d_3_), .A (nx61539z3), .B (
        ENCR_DEV_cnt_init[2]), .C (ENCR_DEV_cnt_init[3])) ;
    AX1 inc_d_5__rename881 (.Y (inc_d_5_), .A (nx61539z2), .B (
        ENCR_DEV_cnt_init[4]), .C (ENCR_DEV_cnt_init[5])) ;
    AX1 inc_d_9__rename882 (.Y (inc_d_9_), .A (nx61539z1), .B (
        ENCR_DEV_cnt_init[8]), .C (ENCR_DEV_cnt_init[9])) ;
    XA1B sclear_and_0_dup_719_rename883 (.Y (sclear_and_0_dup_719), .A (
         ENCR_DEV_err_cnt[0]), .B (ENCR_DEV_prev[2]), .C (ENCR_DEV_prev_6__int)
         ) ;
    XA1C sclear_and_1_dup_720_rename884 (.Y (sclear_and_1_dup_720), .A (
         nx26032z1), .B (ENCR_DEV_err_cnt[1]), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_2_dup_721_rename885 (.Y (sclear_and_2_dup_721), .A (
         ENCR_DEV_err_cnt[2]), .B (nx16750z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_3_dup_722_rename886 (.Y (sclear_and_3_dup_722), .A (nx6004z1
         ), .B (ENCR_DEV_err_cnt[3]), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_4_dup_723_rename887 (.Y (sclear_and_4_dup_723), .A (
         ENCR_DEV_err_cnt[4]), .B (nx36778z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_5_dup_724_rename888 (.Y (sclear_and_5_dup_724), .A (
         ENCR_DEV_err_cnt[5]), .B (nx51512z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_6_dup_725_rename889 (.Y (sclear_and_6_dup_725), .A (
         ENCR_DEV_err_cnt[6]), .B (nx56806z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_7_dup_726_rename890 (.Y (sclear_and_7_dup_726), .A (
         ENCR_DEV_err_cnt[7]), .B (nx31484z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_8_dup_727_rename891 (.Y (sclear_and_8_dup_727), .A (
         ENCR_DEV_err_cnt[8]), .B (nx11298z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_9_dup_728_rename892 (.Y (sclear_and_9_dup_728), .A (
         ENCR_DEV_err_cnt[9]), .B (nx8414z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_10_dup_729_rename893 (.Y (sclear_and_10_dup_729), .A (
         ENCR_DEV_err_cnt[10]), .B (nx5753z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_11_dup_730_rename894 (.Y (sclear_and_11_dup_730), .A (
         ENCR_DEV_err_cnt[11]), .B (nx36042z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_12_dup_731_rename895 (.Y (sclear_and_12_dup_731), .A (
         ENCR_DEV_err_cnt[12]), .B (nx52248z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_13_dup_732_rename896 (.Y (sclear_and_13_dup_732), .A (
         ENCR_DEV_err_cnt[13]), .B (nx56070z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_14_dup_733_rename897 (.Y (sclear_and_14_dup_733), .A (
         ENCR_DEV_err_cnt[14]), .B (nx32220z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_15_dup_734_rename898 (.Y (sclear_and_15_dup_734), .A (
         ENCR_DEV_err_cnt[15]), .B (nx10562z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_16_dup_735_rename899 (.Y (sclear_and_16_dup_735), .A (
         ENCR_DEV_err_cnt[16]), .B (nx12192z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_17_dup_736_rename900 (.Y (sclear_and_17_dup_736), .A (
         ENCR_DEV_err_cnt[17]), .B (nx34946z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_18_dup_737_rename901 (.Y (sclear_and_18_dup_737), .A (
         ENCR_DEV_err_cnt[18]), .B (nx7836z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_19_dup_738_rename902 (.Y (sclear_and_19_dup_738), .A (
         nx14918z1), .B (ENCR_DEV_err_cnt[19]), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_20_dup_739_rename903 (.Y (sclear_and_20_dup_739), .A (
         ENCR_DEV_err_cnt[20]), .B (nx49501z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_21_dup_740_rename904 (.Y (sclear_and_21_dup_740), .A (
         ENCR_DEV_err_cnt[21]), .B (nx39776z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_22_dup_741_rename905 (.Y (sclear_and_22_dup_741), .A (
         ENCR_DEV_err_cnt[22]), .B (nx3006z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_23_dup_742_rename906 (.Y (sclear_and_23_dup_742), .A (
         ENCR_DEV_err_cnt[23]), .B (nx19748z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_24_dup_743_rename907 (.Y (sclear_and_24_dup_743), .A (
         ENCR_DEV_err_cnt[24]), .B (NOT_a_0__dup_3643), .C (ENCR_DEV_prev_6__int
         )) ;
    XA1C sclear_and_25_dup_744_rename908 (.Y (sclear_and_25_dup_744), .A (
         ENCR_DEV_err_cnt[25]), .B (NOT_a_0__dup_3648), .C (ENCR_DEV_prev_6__int
         )) ;
    XA1C sclear_and_26_dup_745_rename909 (.Y (sclear_and_26_dup_745), .A (
         ENCR_DEV_err_cnt[26]), .B (NOT_a_0__dup_3653), .C (ENCR_DEV_prev_6__int
         )) ;
    XA1C sclear_and_27_dup_746_rename910 (.Y (sclear_and_27_dup_746), .A (
         ENCR_DEV_err_cnt[27]), .B (NOT_a_0__dup_3658), .C (ENCR_DEV_prev_6__int
         )) ;
    XA1C sclear_and_28_dup_747_rename911 (.Y (sclear_and_28_dup_747), .A (
         ENCR_DEV_err_cnt[28]), .B (NOT_a_0__dup_3632), .C (ENCR_DEV_prev_6__int
         )) ;
    XA1C sclear_and_29_dup_748_rename912 (.Y (sclear_and_29_dup_748), .A (
         ENCR_DEV_err_cnt[29]), .B (NOT_a_0__dup_3638), .C (ENCR_DEV_prev_6__int
         )) ;
    XA1C sclear_and_30_dup_749_rename913 (.Y (sclear_and_30_dup_749), .A (
         ENCR_DEV_err_cnt[30]), .B (NOT_a_0_), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_31_dup_750_rename914 (.Y (sclear_and_31_dup_750), .A (
         ENCR_DEV_err_cnt[31]), .B (NOT_a_0__dup_3626), .C (ENCR_DEV_prev_6__int
         )) ;
    XA1C sclear_and_32_dup_751_rename915 (.Y (sclear_and_32_dup_751), .A (
         ENCR_DEV_err_cnt[32]), .B (nx7276z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_33_dup_752_rename916 (.Y (sclear_and_33_dup_752), .A (
         ENCR_DEV_err_cnt[33]), .B (nx35506z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_34_dup_753_rename917 (.Y (sclear_and_34_dup_753), .A (
         ENCR_DEV_err_cnt[34]), .B (nx52784z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_35_dup_754_rename918 (.Y (sclear_and_35_dup_754), .A (
         ENCR_DEV_err_cnt[35]), .B (nx55534z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_36_dup_755_rename919 (.Y (sclear_and_36_dup_755), .A (
         ENCR_DEV_err_cnt[36]), .B (nx32756z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_37_dup_756_rename920 (.Y (sclear_and_37_dup_756), .A (
         ENCR_DEV_err_cnt[37]), .B (nx55510z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_38_dup_757_rename921 (.Y (sclear_and_38_dup_757), .A (
         ENCR_DEV_err_cnt[38]), .B (nx52808z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_39_dup_758_rename922 (.Y (sclear_and_39_dup_758), .A (
         ENCR_DEV_err_cnt[39]), .B (nx35482z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_40_dup_759_rename923 (.Y (sclear_and_40_dup_759), .A (
         ENCR_DEV_err_cnt[40]), .B (nx28937z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_41_dup_760_rename924 (.Y (sclear_and_41_dup_760), .A (
         ENCR_DEV_err_cnt[41]), .B (nx60340z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_42_dup_761_rename925 (.Y (sclear_and_42_dup_761), .A (
         ENCR_DEV_err_cnt[42]), .B (nx47978z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_43_dup_762_rename926 (.Y (sclear_and_43_dup_762), .A (
         ENCR_DEV_err_cnt[43]), .B (nx40312z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_44_dup_763_rename927 (.Y (sclear_and_44_dup_763), .A (
         ENCR_DEV_err_cnt[44]), .B (nx2470z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_45_dup_764_rename928 (.Y (sclear_and_45_dup_764), .A (
         ENCR_DEV_err_cnt[45]), .B (nx20284z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_46_dup_765_rename929 (.Y (sclear_and_46_dup_765), .A (
         ENCR_DEV_err_cnt[46]), .B (nx22498z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_47_dup_766_rename930 (.Y (sclear_and_47_dup_766), .A (
         ENCR_DEV_err_cnt[47]), .B (nx65280z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_48_dup_767_rename931 (.Y (sclear_and_48_dup_767), .A (
         ENCR_DEV_err_cnt[48]), .B (nx23010z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_49_dup_768_rename932 (.Y (sclear_and_49_dup_768), .A (
         ENCR_DEV_err_cnt[49]), .B (nx19772z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_50_dup_769_rename933 (.Y (sclear_and_50_dup_769), .A (
         ENCR_DEV_err_cnt[50]), .B (nx46881z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_51_dup_770_rename934 (.Y (sclear_and_51_dup_770), .A (
         nx60450z1), .B (ENCR_DEV_err_cnt[51]), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_52_dup_771_rename935 (.Y (sclear_and_52_dup_771), .A (
         ENCR_DEV_err_cnt[52]), .B (nx27840z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_53_dup_772_rename936 (.Y (sclear_and_53_dup_772), .A (
         ENCR_DEV_err_cnt[53]), .B (nx14942z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_54_dup_773_rename937 (.Y (sclear_and_54_dup_773), .A (
         ENCR_DEV_err_cnt[54]), .B (nx7812z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_55_dup_774_rename938 (.Y (sclear_and_55_dup_774), .A (
         ENCR_DEV_err_cnt[55]), .B (nx34970z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_56_dup_775_rename939 (.Y (sclear_and_56_dup_775), .A (
         ENCR_DEV_err_cnt[56]), .B (nx12216z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_57_dup_776_rename940 (.Y (sclear_and_57_dup_776), .A (
         ENCR_DEV_err_cnt[57]), .B (nx10538z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_58_dup_777_rename941 (.Y (sclear_and_58_dup_777), .A (
         ENCR_DEV_err_cnt[58]), .B (nx32244z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_59_dup_778_rename942 (.Y (sclear_and_59_dup_778), .A (
         ENCR_DEV_err_cnt[59]), .B (nx56046z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_60_dup_779_rename943 (.Y (sclear_and_60_dup_779), .A (
         ENCR_DEV_err_cnt[60]), .B (nx8373z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_61_dup_780_rename944 (.Y (sclear_and_61_dup_780), .A (
         ENCR_DEV_err_cnt[61]), .B (nx15368z1), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_62_dup_781_rename945 (.Y (sclear_and_62_dup_781), .A (
         nx27414z1), .B (ENCR_DEV_err_cnt[62]), .C (ENCR_DEV_prev_6__int)) ;
    XA1C sclear_and_63_dup_782_rename946 (.Y (sclear_and_63_dup_782), .A (
         nx60876z1), .B (ENCR_DEV_err_cnt[63]), .C (ENCR_DEV_prev_6__int)) ;
    NAND2 NOT_ix26032z24338 (.Y (nx26032z1), .A (ENCR_DEV_prev[2]), .B (
          ENCR_DEV_err_cnt[0])) ;
    NAND3 NOT_ix16750z24337 (.Y (nx16750z1), .A (ENCR_DEV_prev[2]), .B (
          ENCR_DEV_err_cnt[0]), .C (ENCR_DEV_err_cnt[1])) ;
    NAND2 NOT_ix8414z24340 (.Y (nx8414z3), .A (ENCR_DEV_err_cnt[2]), .B (
          ENCR_DEV_err_cnt[1])) ;
    NAND2 NOT_a_10__rename947 (.Y (NOT_a_10_), .A (ENCR_DEV_err_cnt[3]), .B (
          ENCR_DEV_err_cnt[2])) ;
    NAND2 NOT_ix8414z24341 (.Y (nx8414z4), .A (ENCR_DEV_err_cnt[4]), .B (
          ENCR_DEV_err_cnt[3])) ;
    NAND2 NOT_ix11298z24339 (.Y (nx11298z2), .A (ENCR_DEV_err_cnt[5]), .B (
          ENCR_DEV_err_cnt[4])) ;
    NAND2 NOT_ix11298z24340 (.Y (nx11298z3), .A (ENCR_DEV_err_cnt[7]), .B (
          ENCR_DEV_err_cnt[6])) ;
    NAND2 NOT_ix8414z24343 (.Y (nx8414z6), .A (ENCR_DEV_err_cnt[8]), .B (
          ENCR_DEV_err_cnt[7])) ;
    NAND2 NOT_ix49501z24342 (.Y (nx49501z4), .A (ENCR_DEV_err_cnt[9]), .B (
          ENCR_DEV_err_cnt[8])) ;
    NAND2 NOT_ix56070z24340 (.Y (nx56070z3), .A (ENCR_DEV_err_cnt[12]), .B (
          ENCR_DEV_err_cnt[11])) ;
    NAND2 NOT_ix49501z24345 (.Y (nx49501z7), .A (ENCR_DEV_err_cnt[13]), .B (
          ENCR_DEV_err_cnt[12])) ;
    NAND2 NOT_ix34946z24342 (.Y (nx34946z4), .A (ENCR_DEV_err_cnt[16]), .B (
          ENCR_DEV_err_cnt[15])) ;
    NAND2 NOT_ix49501z24347 (.Y (nx49501z9), .A (ENCR_DEV_err_cnt[17]), .B (
          ENCR_DEV_err_cnt[16])) ;
    NAND2 NOT_ix8414z24346 (.Y (nx8414z9), .A (ENCR_DEV_err_cnt[20]), .B (
          ENCR_DEV_err_cnt[19])) ;
    NAND2 NOT_ix8409z24342 (.Y (nx8409z4), .A (ENCR_DEV_err_cnt[21]), .B (
          ENCR_DEV_err_cnt[20])) ;
    NAND2 NOT_ix8414z24348 (.Y (nx8414z11), .A (ENCR_DEV_err_cnt[24]), .B (
          ENCR_DEV_err_cnt[23])) ;
    NAND2 NOT_ix11504z24343 (.Y (nx11504z5), .A (ENCR_DEV_err_cnt[25]), .B (
          ENCR_DEV_err_cnt[24])) ;
    NAND2 NOT_ix7417z24340 (.Y (nx7417z3), .A (ENCR_DEV_err_cnt[28]), .B (
          ENCR_DEV_err_cnt[27])) ;
    NAND2 NOT_ix11504z24345 (.Y (nx11504z7), .A (ENCR_DEV_err_cnt[29]), .B (
          ENCR_DEV_err_cnt[28])) ;
    NAND2 NOT_ix35506z24344 (.Y (nx35506z6), .A (ENCR_DEV_err_cnt[32]), .B (
          ENCR_DEV_err_cnt[31])) ;
    NAND2 NOT_ix11504z24351 (.Y (nx11504z13), .A (ENCR_DEV_err_cnt[33]), .B (
          ENCR_DEV_err_cnt[32])) ;
    NAND2 NOT_ix55510z24342 (.Y (nx55510z4), .A (ENCR_DEV_err_cnt[36]), .B (
          ENCR_DEV_err_cnt[35])) ;
    NAND2 NOT_ix11504z24353 (.Y (nx11504z15), .A (ENCR_DEV_err_cnt[37]), .B (
          ENCR_DEV_err_cnt[36])) ;
    NAND2 NOT_ix40554z24340 (.Y (nx40554z3), .A (ENCR_DEV_err_cnt[40]), .B (
          ENCR_DEV_err_cnt[39])) ;
    NAND2 NOT_ix41545z24339 (.Y (nx41545z2), .A (ENCR_DEV_err_cnt[41]), .B (
          ENCR_DEV_err_cnt[40])) ;
    NAND2 NOT_ix20284z24343 (.Y (nx20284z5), .A (ENCR_DEV_err_cnt[44]), .B (
          ENCR_DEV_err_cnt[43])) ;
    NAND2 NOT_ix41545z24341 (.Y (nx41545z4), .A (ENCR_DEV_err_cnt[45]), .B (
          ENCR_DEV_err_cnt[44])) ;
    NAND2 NOT_ix19772z24342 (.Y (nx19772z4), .A (ENCR_DEV_err_cnt[48]), .B (
          ENCR_DEV_err_cnt[47])) ;
    NAND2 NOT_ix7423z24338 (.Y (nx7423z1), .A (ENCR_DEV_err_cnt[49]), .B (
          ENCR_DEV_err_cnt[48])) ;
    NAND2 NOT_ix7418z24338 (.Y (nx7418z1), .A (ENCR_DEV_err_cnt[52]), .B (
          ENCR_DEV_err_cnt[51])) ;
    NAND2 NOT_ix9408z24338 (.Y (nx9408z1), .A (ENCR_DEV_err_cnt[53]), .B (
          ENCR_DEV_err_cnt[52])) ;
    NAND2 NOT_ix8415z24338 (.Y (nx8415z1), .A (ENCR_DEV_err_cnt[56]), .B (
          ENCR_DEV_err_cnt[55])) ;
    NAND2 NOT_a_4__dup_3628_rename948 (.Y (NOT_a_4__dup_3628), .A (
          ENCR_DEV_err_cnt[57]), .B (ENCR_DEV_err_cnt[56])) ;
    NAND2 NOT_a_4__rename949 (.Y (NOT_a_4_), .A (ENCR_DEV_err_cnt[59]), .B (
          ENCR_DEV_err_cnt[58])) ;
    NAND2 NOT_a_4__dup_3622_rename950 (.Y (NOT_a_4__dup_3622), .A (
          ENCR_DEV_err_cnt[60]), .B (ENCR_DEV_err_cnt[59])) ;
    NAND3A NOT_ix6004z50930 (.Y (nx6004z1), .A (nx26032z1), .B (
           ENCR_DEV_err_cnt[2]), .C (ENCR_DEV_err_cnt[1])) ;
    NAND3A NOT_ix36778z50930 (.Y (nx36778z1), .A (nx16750z1), .B (
           ENCR_DEV_err_cnt[3]), .C (ENCR_DEV_err_cnt[2])) ;
    NAND3A NOT_ix31484z50931 (.Y (nx31484z2), .A (nx8414z4), .B (
           ENCR_DEV_err_cnt[6]), .C (ENCR_DEV_err_cnt[5])) ;
    NAND3A NOT_a_9__rename951 (.Y (NOT_a_9_), .A (nx11298z2), .B (
           ENCR_DEV_err_cnt[7]), .C (ENCR_DEV_err_cnt[6])) ;
    NAND3A NOT_ix8414z50934 (.Y (nx8414z5), .A (nx8414z6), .B (
           ENCR_DEV_err_cnt[5]), .C (ENCR_DEV_err_cnt[6])) ;
    NAND3A NOT_ix5753z50932 (.Y (nx5753z3), .A (nx11298z3), .B (
           ENCR_DEV_err_cnt[8]), .C (ENCR_DEV_err_cnt[9])) ;
    NAND3A NOT_ix36042z50931 (.Y (nx36042z2), .A (nx8414z6), .B (
           ENCR_DEV_err_cnt[10]), .C (ENCR_DEV_err_cnt[9])) ;
    NAND3A NOT_ix49501z50937 (.Y (nx49501z3), .A (nx49501z4), .B (
           ENCR_DEV_err_cnt[11]), .C (ENCR_DEV_err_cnt[10])) ;
    NAND3A NOT_ix56070z50931 (.Y (nx56070z2), .A (nx56070z3), .B (
           ENCR_DEV_err_cnt[9]), .C (ENCR_DEV_err_cnt[10])) ;
    NAND3A NOT_ix32220z50931 (.Y (nx32220z2), .A (nx49501z7), .B (
           ENCR_DEV_err_cnt[10]), .C (ENCR_DEV_err_cnt[11])) ;
    NAND3A NOT_ix10562z50932 (.Y (nx10562z3), .A (nx56070z3), .B (
           ENCR_DEV_err_cnt[14]), .C (ENCR_DEV_err_cnt[13])) ;
    NAND3A NOT_ix49501z50936 (.Y (nx49501z6), .A (nx49501z7), .B (
           ENCR_DEV_err_cnt[15]), .C (ENCR_DEV_err_cnt[14])) ;
    NAND3A NOT_ix34946z50937 (.Y (nx34946z3), .A (nx34946z4), .B (
           ENCR_DEV_err_cnt[14]), .C (ENCR_DEV_err_cnt[13])) ;
    NAND3A NOT_ix7836z50937 (.Y (nx7836z3), .A (nx49501z9), .B (
           ENCR_DEV_err_cnt[14]), .C (ENCR_DEV_err_cnt[15])) ;
    NAND3A NOT_ix14918z50939 (.Y (nx14918z4), .A (nx34946z4), .B (
           ENCR_DEV_err_cnt[18]), .C (ENCR_DEV_err_cnt[17])) ;
    NAND3A NOT_ix49501z50938 (.Y (nx49501z8), .A (nx49501z9), .B (
           ENCR_DEV_err_cnt[19]), .C (ENCR_DEV_err_cnt[18])) ;
    NAND3A NOT_ix8414z50937 (.Y (nx8414z8), .A (nx8414z9), .B (
           ENCR_DEV_err_cnt[17]), .C (ENCR_DEV_err_cnt[18])) ;
    NAND3A NOT_ix3006z50939 (.Y (nx3006z4), .A (nx8409z4), .B (
           ENCR_DEV_err_cnt[18]), .C (ENCR_DEV_err_cnt[19])) ;
    NAND3A NOT_ix19748z50937 (.Y (nx19748z3), .A (nx8414z9), .B (
           ENCR_DEV_err_cnt[22]), .C (ENCR_DEV_err_cnt[21])) ;
    NAND3A NOT_ix8409z50937 (.Y (nx8409z3), .A (nx8409z4), .B (
           ENCR_DEV_err_cnt[23]), .C (ENCR_DEV_err_cnt[22])) ;
    NAND3A NOT_ix8414z50939 (.Y (nx8414z10), .A (nx8414z11), .B (
           ENCR_DEV_err_cnt[21]), .C (ENCR_DEV_err_cnt[22])) ;
    NAND3A NOT_ix9406z50931 (.Y (nx9406z2), .A (nx11504z5), .B (
           ENCR_DEV_err_cnt[23]), .C (ENCR_DEV_err_cnt[22])) ;
    NAND3A NOT_ix9411z50931 (.Y (nx9411z2), .A (nx8414z11), .B (
           ENCR_DEV_err_cnt[26]), .C (ENCR_DEV_err_cnt[25])) ;
    NAND3A NOT_ix11504z50934 (.Y (nx11504z4), .A (nx11504z5), .B (
           ENCR_DEV_err_cnt[27]), .C (ENCR_DEV_err_cnt[26])) ;
    NAND3A NOT_ix7417z50931 (.Y (nx7417z2), .A (nx7417z3), .B (
           ENCR_DEV_err_cnt[25]), .C (ENCR_DEV_err_cnt[26])) ;
    NAND3A NOT_ix32078z50931 (.Y (nx32078z2), .A (nx11504z7), .B (
           ENCR_DEV_err_cnt[27]), .C (ENCR_DEV_err_cnt[26])) ;
    NAND3A NOT_ix6418z50932 (.Y (nx6418z3), .A (nx7417z3), .B (
           ENCR_DEV_err_cnt[30]), .C (ENCR_DEV_err_cnt[29])) ;
    NAND3A NOT_ix11504z50936 (.Y (nx11504z6), .A (nx11504z7), .B (
           ENCR_DEV_err_cnt[31]), .C (ENCR_DEV_err_cnt[30])) ;
    NAND3A NOT_ix35506z50941 (.Y (nx35506z5), .A (nx35506z6), .B (
           ENCR_DEV_err_cnt[29]), .C (ENCR_DEV_err_cnt[30])) ;
    NAND3A NOT_ix52784z50941 (.Y (nx52784z5), .A (nx11504z13), .B (
           ENCR_DEV_err_cnt[31]), .C (ENCR_DEV_err_cnt[30])) ;
    NAND3A NOT_ix55534z50939 (.Y (nx55534z4), .A (nx35506z6), .B (
           ENCR_DEV_err_cnt[34]), .C (ENCR_DEV_err_cnt[33])) ;
    NAND3A NOT_ix11504z50942 (.Y (nx11504z12), .A (nx11504z13), .B (
           ENCR_DEV_err_cnt[35]), .C (ENCR_DEV_err_cnt[34])) ;
    NAND3A NOT_ix55510z50937 (.Y (nx55510z3), .A (nx55510z4), .B (
           ENCR_DEV_err_cnt[33]), .C (ENCR_DEV_err_cnt[34])) ;
    NAND3A NOT_ix52808z50937 (.Y (nx52808z3), .A (nx11504z15), .B (
           ENCR_DEV_err_cnt[34]), .C (ENCR_DEV_err_cnt[35])) ;
    NAND3A NOT_ix35482z50937 (.Y (nx35482z3), .A (nx55510z4), .B (
           ENCR_DEV_err_cnt[38]), .C (ENCR_DEV_err_cnt[37])) ;
    NAND3A NOT_ix11504z50944 (.Y (nx11504z14), .A (nx11504z15), .B (
           ENCR_DEV_err_cnt[39]), .C (ENCR_DEV_err_cnt[38])) ;
    NAND3A NOT_ix40554z50931 (.Y (nx40554z2), .A (nx40554z3), .B (
           ENCR_DEV_err_cnt[37]), .C (ENCR_DEV_err_cnt[38])) ;
    NAND3A NOT_ix39562z50931 (.Y (nx39562z2), .A (nx41545z2), .B (
           ENCR_DEV_err_cnt[38]), .C (ENCR_DEV_err_cnt[39])) ;
    NAND3A NOT_ix39557z50931 (.Y (nx39557z2), .A (nx40554z3), .B (
           ENCR_DEV_err_cnt[42]), .C (ENCR_DEV_err_cnt[41])) ;
    NAND3A NOT_ix41545z50930 (.Y (nx41545z1), .A (nx41545z2), .B (
           ENCR_DEV_err_cnt[43]), .C (ENCR_DEV_err_cnt[42])) ;
    NAND3A NOT_ix20284z50934 (.Y (nx20284z4), .A (nx20284z5), .B (
           ENCR_DEV_err_cnt[41]), .C (ENCR_DEV_err_cnt[42])) ;
    NAND3A NOT_ix22498z50934 (.Y (nx22498z4), .A (nx41545z4), .B (
           ENCR_DEV_err_cnt[42]), .C (ENCR_DEV_err_cnt[43])) ;
    NAND3A NOT_ix65280z50933 (.Y (nx65280z3), .A (nx20284z5), .B (
           ENCR_DEV_err_cnt[46]), .C (ENCR_DEV_err_cnt[45])) ;
    NAND3A NOT_ix41545z50932 (.Y (nx41545z3), .A (nx41545z4), .B (
           ENCR_DEV_err_cnt[47]), .C (ENCR_DEV_err_cnt[46])) ;
    NAND3A NOT_ix19772z50937 (.Y (nx19772z3), .A (nx19772z4), .B (
           ENCR_DEV_err_cnt[45]), .C (ENCR_DEV_err_cnt[46])) ;
    NAND3A NOT_ix42542z50930 (.Y (nx42542z1), .A (nx7423z1), .B (
           ENCR_DEV_err_cnt[47]), .C (ENCR_DEV_err_cnt[46])) ;
    NAND3A NOT_ix60450z50937 (.Y (nx60450z3), .A (nx19772z4), .B (
           ENCR_DEV_err_cnt[50]), .C (ENCR_DEV_err_cnt[49])) ;
    NAND3A NOT_a_3__dup_3640_rename952 (.Y (NOT_a_3__dup_3640), .A (nx7423z1), .B (
           ENCR_DEV_err_cnt[51]), .C (ENCR_DEV_err_cnt[50])) ;
    NAND3A NOT_a_3__dup_3645_rename953 (.Y (NOT_a_3__dup_3645), .A (nx7418z1), .B (
           ENCR_DEV_err_cnt[49]), .C (ENCR_DEV_err_cnt[50])) ;
    NAND3A NOT_a_3__dup_3650_rename954 (.Y (NOT_a_3__dup_3650), .A (nx9408z1), .B (
           ENCR_DEV_err_cnt[51]), .C (ENCR_DEV_err_cnt[50])) ;
    NAND3A NOT_a_3__dup_3655_rename955 (.Y (NOT_a_3__dup_3655), .A (nx7418z1), .B (
           ENCR_DEV_err_cnt[54]), .C (ENCR_DEV_err_cnt[53])) ;
    NAND3A NOT_a_3__dup_3629_rename956 (.Y (NOT_a_3__dup_3629), .A (nx9408z1), .B (
           ENCR_DEV_err_cnt[55]), .C (ENCR_DEV_err_cnt[54])) ;
    NAND3A NOT_a_3__dup_3635_rename957 (.Y (NOT_a_3__dup_3635), .A (nx8415z1), .B (
           ENCR_DEV_err_cnt[53]), .C (ENCR_DEV_err_cnt[54])) ;
    NAND3A NOT_a_3__rename958 (.Y (NOT_a_3_), .A (NOT_a_4__dup_3628), .B (
           ENCR_DEV_err_cnt[55]), .C (ENCR_DEV_err_cnt[54])) ;
    NAND3A NOT_a_3__dup_3623_rename959 (.Y (NOT_a_3__dup_3623), .A (nx8415z1), .B (
           ENCR_DEV_err_cnt[58]), .C (ENCR_DEV_err_cnt[57])) ;
    NAND3C NOT_ix51512z50932 (.Y (nx51512z1), .A (nx26032z1), .B (nx8414z3), .C (
           nx8414z4)) ;
    NAND3C NOT_ix56806z50932 (.Y (nx56806z1), .A (nx16750z1), .B (NOT_a_10_), .C (
           nx11298z2)) ;
    NAND2B NOT_ix31484z49934 (.Y (nx31484z1), .A (nx6004z1), .B (nx31484z2)) ;
    NAND3C NOT_ix11298z50932 (.Y (nx11298z1), .A (nx11298z2), .B (nx11298z3), .C (
           nx36778z1)) ;
    NAND3C NOT_ix8414z50933 (.Y (nx8414z2), .A (nx8414z3), .B (nx8414z4), .C (
           nx8414z5)) ;
    NAND3C NOT_ix5753z50933 (.Y (nx5753z2), .A (NOT_a_10_), .B (nx11298z2), .C (
           nx5753z3)) ;
    NAND2B NOT_ix10562z49935 (.Y (nx10562z2), .A (nx36042z2), .B (nx10562z3)) ;
    NAND2B NOT_ix34946z49935 (.Y (nx34946z2), .A (nx56070z2), .B (nx34946z3)) ;
    NAND2B NOT_ix7836z49935 (.Y (nx7836z2), .A (nx7836z3), .B (nx32220z2)) ;
    NAND2B NOT_ix14918z49936 (.Y (nx14918z3), .A (nx10562z3), .B (nx14918z4)) ;
    NAND2B NOT_ix49501z49939 (.Y (nx49501z5), .A (nx49501z6), .B (nx49501z8)) ;
    NAND2B NOT_ix39776z49936 (.Y (nx39776z3), .A (nx34946z3), .B (nx8414z8)) ;
    NAND2B NOT_ix3006z49936 (.Y (nx3006z3), .A (nx7836z3), .B (nx3006z4)) ;
    NAND2B NOT_ix8409z49935 (.Y (nx8409z2), .A (nx49501z8), .B (nx8409z3)) ;
    NAND2B NOT_ix7411z49934 (.Y (nx7411z1), .A (nx8409z3), .B (nx11504z4)) ;
    NAND2B NOT_ix7417z49934 (.Y (nx7417z1), .A (nx8414z10), .B (nx7417z2)) ;
    NAND2B NOT_ix32078z49934 (.Y (nx32078z1), .A (nx9406z2), .B (nx32078z2)) ;
    NAND2B NOT_ix6418z49935 (.Y (nx6418z2), .A (nx9411z2), .B (nx6418z3)) ;
    NAND2B NOT_ix11504z49937 (.Y (nx11504z3), .A (nx11504z4), .B (nx11504z6)) ;
    NAND2B NOT_ix35506z49937 (.Y (nx35506z4), .A (nx35506z5), .B (nx7417z2)) ;
    NAND2B NOT_ix52784z49937 (.Y (nx52784z4), .A (nx32078z2), .B (nx52784z5)) ;
    NAND2B NOT_ix55534z49936 (.Y (nx55534z3), .A (nx6418z3), .B (nx55534z4)) ;
    NAND2B NOT_ix41557z49934 (.Y (nx41557z1), .A (nx11504z6), .B (nx11504z12)) ;
    NAND2B NOT_ix11504z49945 (.Y (nx11504z11), .A (nx11504z12), .B (nx11504z14)
           ) ;
    NAND2B NOT_ix40554z49934 (.Y (nx40554z1), .A (nx55510z3), .B (nx40554z2)) ;
    NAND2B NOT_ix39562z49934 (.Y (nx39562z1), .A (nx52808z3), .B (nx39562z2)) ;
    NAND2B NOT_ix39557z49934 (.Y (nx39557z1), .A (nx35482z3), .B (nx39557z2)) ;
    NAND2B NOT_ix20284z49937 (.Y (nx20284z3), .A (nx40554z2), .B (nx20284z4)) ;
    NAND2B NOT_ix22498z49937 (.Y (nx22498z3), .A (nx39562z2), .B (nx22498z4)) ;
    NAND2B NOT_ix65280z49936 (.Y (nx65280z2), .A (nx39557z2), .B (nx65280z3)) ;
    NAND2B NOT_a_2__dup_3641_rename960 (.Y (NOT_a_2__dup_3641), .A (nx41545z1), 
           .B (nx41545z3)) ;
    NAND2B NOT_a_2__dup_3646_rename961 (.Y (NOT_a_2__dup_3646), .A (nx19772z3), 
           .B (nx20284z4)) ;
    NAND2B NOT_a_2__dup_3651_rename962 (.Y (NOT_a_2__dup_3651), .A (nx22498z4), 
           .B (nx42542z1)) ;
    NAND2B NOT_a_2__dup_3656_rename963 (.Y (NOT_a_2__dup_3656), .A (nx65280z3), 
           .B (nx60450z3)) ;
    NAND2B NOT_a_2__dup_3630_rename964 (.Y (NOT_a_2__dup_3630), .A (nx41545z3), 
           .B (NOT_a_3__dup_3640)) ;
    NAND2B NOT_a_2__dup_3636_rename965 (.Y (NOT_a_2__dup_3636), .A (nx19772z3), 
           .B (NOT_a_3__dup_3645)) ;
    NAND2B NOT_a_2__rename966 (.Y (NOT_a_2_), .A (nx42542z1), .B (
           NOT_a_3__dup_3650)) ;
    NAND2B NOT_a_2__dup_3624_rename967 (.Y (NOT_a_2__dup_3624), .A (nx60450z3), 
           .B (NOT_a_3__dup_3655)) ;
    NAND3A NOT_ix8414z50930 (.Y (nx8414z1), .A (nx8414z2), .B (
           ENCR_DEV_err_cnt[0]), .C (ENCR_DEV_prev[2])) ;
    NAND3B NOT_ix5753z50931 (.Y (nx5753z1), .A (nx26032z1), .B (nx5753z2), .C (
           ENCR_DEV_err_cnt[1])) ;
    NAND3C NOT_ix36042z50932 (.Y (nx36042z1), .A (nx31484z2), .B (nx36042z2), .C (
           nx6004z1)) ;
    NAND3C NOT_ix52248z50932 (.Y (nx52248z1), .A (nx36778z1), .B (NOT_a_9_), .C (
           nx49501z3)) ;
    NAND3C NOT_ix56070z50932 (.Y (nx56070z1), .A (nx51512z1), .B (nx8414z5), .C (
           nx56070z2)) ;
    NAND3C NOT_ix32220z50932 (.Y (nx32220z1), .A (nx56806z1), .B (nx5753z3), .C (
           nx32220z2)) ;
    NAND3C NOT_ix12192z50932 (.Y (nx12192z1), .A (nx11298z1), .B (nx49501z3), .C (
           nx49501z6)) ;
    NAND3C NOT_ix35506z50933 (.Y (nx35506z2), .A (nx8414z2), .B (nx56070z2), .C (
           nx34946z3)) ;
    NAND3C NOT_ix52784z50933 (.Y (nx52784z2), .A (nx5753z2), .B (nx32220z2), .C (
           nx7836z3)) ;
    NAND3C NOT_ix14918z50933 (.Y (nx14918z2), .A (nx31484z2), .B (nx36042z2), .C (
           nx14918z3)) ;
    NAND3C NOT_ix49501z50933 (.Y (nx49501z2), .A (NOT_a_9_), .B (nx49501z3), .C (
           nx49501z5)) ;
    NAND3C NOT_ix39776z50933 (.Y (nx39776z2), .A (nx8414z5), .B (nx56070z2), .C (
           nx39776z3)) ;
    NAND3C NOT_ix3006z50933 (.Y (nx3006z2), .A (nx3006z3), .B (nx5753z3), .C (
           nx32220z2)) ;
    NAND3C NOT_ix19748z50933 (.Y (nx19748z2), .A (nx14918z4), .B (nx19748z3), .C (
           nx10562z2)) ;
    NAND3C NOT_ix8409z50932 (.Y (nx8409z1), .A (nx49501z3), .B (nx49501z6), .C (
           nx8409z2)) ;
    NAND3C NOT_ix8414z50938 (.Y (nx8414z7), .A (nx8414z8), .B (nx8414z10), .C (
           nx34946z2)) ;
    NAND3C NOT_ix9406z50932 (.Y (nx9406z1), .A (nx3006z4), .B (nx9406z2), .C (
           nx7836z2)) ;
    NAND3C NOT_ix9411z50932 (.Y (nx9411z1), .A (nx14918z3), .B (nx19748z3), .C (
           nx9411z2)) ;
    NAND3C NOT_ix2470z50933 (.Y (nx2470z2), .A (nx49501z5), .B (nx8409z3), .C (
           nx11504z4)) ;
    NAND3C NOT_ix35506z50934 (.Y (nx35506z3), .A (nx8414z8), .B (nx8414z10), .C (
           nx35506z4)) ;
    NAND3C NOT_ix52784z50934 (.Y (nx52784z3), .A (nx3006z4), .B (nx9406z2), .C (
           nx52784z4)) ;
    NAND3C NOT_ix55534z50933 (.Y (nx55534z2), .A (nx19748z3), .B (nx9411z2), .C (
           nx55534z3)) ;
    NAND3C NOT_ix32756z50933 (.Y (nx32756z2), .A (nx11504z6), .B (nx11504z12), .C (
           nx7411z1)) ;
    NAND3C NOT_ix55510z50933 (.Y (nx55510z2), .A (nx35506z5), .B (nx55510z3), .C (
           nx7417z1)) ;
    NAND3C NOT_ix52808z50933 (.Y (nx52808z2), .A (nx32078z1), .B (nx52784z5), .C (
           nx52808z3)) ;
    NAND3C NOT_ix35482z50933 (.Y (nx35482z2), .A (nx55534z4), .B (nx35482z3), .C (
           nx6418z2)) ;
    NAND3C NOT_a_1__dup_3642_rename968 (.Y (NOT_a_1__dup_3642), .A (nx11504z12)
           , .B (nx11504z14), .C (nx11504z3)) ;
    NAND3C NOT_a_1__dup_3647_rename969 (.Y (NOT_a_1__dup_3647), .A (nx35506z5), 
           .B (nx7417z2), .C (nx40554z1)) ;
    NAND3C NOT_a_1__dup_3652_rename970 (.Y (NOT_a_1__dup_3652), .A (nx32078z2), 
           .B (nx52784z5), .C (nx39562z1)) ;
    NAND3C NOT_a_1__dup_3657_rename971 (.Y (NOT_a_1__dup_3657), .A (nx6418z3), .B (
           nx55534z4), .C (nx39557z1)) ;
    NAND3C NOT_a_1__dup_3631_rename972 (.Y (NOT_a_1__dup_3631), .A (nx41557z1), 
           .B (nx11504z14), .C (nx41545z1)) ;
    NAND3C NOT_ix19772z50933 (.Y (nx19772z2), .A (nx40554z1), .B (nx20284z4), .C (
           nx19772z3)) ;
    NAND3C NOT_ix46881z50933 (.Y (nx46881z2), .A (nx52808z3), .B (nx39562z2), .C (
           NOT_a_2__dup_3651)) ;
    NAND3C NOT_ix60450z50933 (.Y (nx60450z2), .A (nx39557z1), .B (nx65280z3), .C (
           nx60450z3)) ;
    NAND3C NOT_ix27840z50933 (.Y (nx27840z2), .A (nx11504z14), .B (nx41545z1), .C (
           NOT_a_2__dup_3630)) ;
    NAND3C NOT_ix14942z50933 (.Y (nx14942z2), .A (NOT_a_2__dup_3636), .B (
           nx40554z2), .C (nx20284z4)) ;
    NAND3C NOT_ix7812z50933 (.Y (nx7812z2), .A (nx39562z2), .B (nx22498z4), .C (
           NOT_a_2_)) ;
    NAND3C NOT_ix34970z50933 (.Y (nx34970z2), .A (nx65280z3), .B (nx39557z2), .C (
           NOT_a_2__dup_3624)) ;
    NAND3C NOT_ix34946z50932 (.Y (nx34946z1), .A (nx26032z1), .B (nx8414z2), .C (
           nx34946z2)) ;
    NAND3C NOT_ix7836z50932 (.Y (nx7836z1), .A (nx5753z2), .B (nx7836z2), .C (
           nx16750z1)) ;
    NAND2B NOT_ix14918z49934 (.Y (nx14918z1), .A (nx6004z1), .B (nx14918z2)) ;
    NAND3C NOT_ix49501z50932 (.Y (nx49501z1), .A (nx16750z1), .B (NOT_a_10_), .C (
           nx49501z2)) ;
    NAND2B NOT_ix39776z49934 (.Y (nx39776z1), .A (nx51512z1), .B (nx39776z2)) ;
    NAND2B NOT_ix3006z49934 (.Y (nx3006z1), .A (nx56806z1), .B (nx3006z2)) ;
    NAND3C NOT_ix19748z50932 (.Y (nx19748z1), .A (nx31484z2), .B (nx6004z1), .C (
           nx19748z2)) ;
    NAND2B NOT_a_0__dup_3643_rename973 (.Y (NOT_a_0__dup_3643), .A (nx11298z1), 
           .B (nx8409z1)) ;
    NAND2B NOT_a_0__dup_3648_rename974 (.Y (NOT_a_0__dup_3648), .A (nx8414z1), .B (
           nx8414z7)) ;
    NAND2B NOT_a_0__dup_3653_rename975 (.Y (NOT_a_0__dup_3653), .A (nx5753z1), .B (
           nx9406z1)) ;
    NAND2B NOT_a_0__dup_3658_rename976 (.Y (NOT_a_0__dup_3658), .A (nx36042z1), 
           .B (nx9411z1)) ;
    NAND3C NOT_a_0__dup_3632_rename977 (.Y (NOT_a_0__dup_3632), .A (nx52248z1), 
           .B (nx49501z5), .C (nx7411z1)) ;
    NAND3C NOT_a_0__dup_3638_rename978 (.Y (NOT_a_0__dup_3638), .A (nx56070z1), 
           .B (nx39776z3), .C (nx7417z1)) ;
    NAND3C NOT_a_0__rename979 (.Y (NOT_a_0_), .A (nx3006z3), .B (nx32078z1), .C (
           nx32220z1)) ;
    NAND2B NOT_a_0__dup_3626_rename980 (.Y (NOT_a_0__dup_3626), .A (nx10562z1), 
           .B (nx6418z1)) ;
    NAND3C NOT_ix7276z50932 (.Y (nx7276z1), .A (nx12192z1), .B (nx8409z2), .C (
           nx11504z3)) ;
    NAND3C NOT_ix20284z50933 (.Y (nx20284z2), .A (nx39776z3), .B (nx7417z1), .C (
           NOT_a_1__dup_3637)) ;
    NAND3C NOT_ix22498z50933 (.Y (nx22498z2), .A (nx3006z3), .B (nx32078z1), .C (
           NOT_a_1_)) ;
    NAND3C NOT_ix23010z50933 (.Y (nx23010z2), .A (NOT_a_7_), .B (nx11504z11), .C (
           NOT_a_2__dup_3641)) ;
    NAND3C NOT_ix35506z50932 (.Y (nx35506z1), .A (nx26032z1), .B (nx35506z2), .C (
           nx35506z3)) ;
    NAND3C NOT_ix52784z50932 (.Y (nx52784z1), .A (nx52784z2), .B (nx16750z1), .C (
           nx52784z3)) ;
    NAND3C NOT_ix55534z50932 (.Y (nx55534z1), .A (nx6004z1), .B (nx14918z2), .C (
           nx55534z2)) ;
    NAND3C NOT_ix32756z50932 (.Y (nx32756z1), .A (nx36778z1), .B (nx49501z2), .C (
           nx32756z2)) ;
    NAND3C NOT_ix55510z50932 (.Y (nx55510z1), .A (nx51512z1), .B (nx39776z2), .C (
           nx55510z2)) ;
    NAND3C NOT_ix52808z50932 (.Y (nx52808z1), .A (nx56806z1), .B (nx3006z2), .C (
           nx52808z2)) ;
    NAND3C NOT_ix35482z50932 (.Y (nx35482z1), .A (nx31484z1), .B (nx19748z2), .C (
           nx35482z2)) ;
    NAND3C NOT_ix28937z50932 (.Y (nx28937z1), .A (nx11298z1), .B (nx8409z1), .C (
           NOT_a_1__dup_3642)) ;
    NAND3C NOT_ix60340z50932 (.Y (nx60340z1), .A (nx8414z7), .B (
           NOT_a_1__dup_3647), .C (nx8414z1)) ;
    NAND3C NOT_ix47978z50932 (.Y (nx47978z1), .A (nx9406z1), .B (
           NOT_a_1__dup_3652), .C (nx5753z1)) ;
    NAND3C NOT_ix40312z50932 (.Y (nx40312z1), .A (nx9411z1), .B (
           NOT_a_1__dup_3657), .C (nx36042z1)) ;
    NAND3C NOT_ix2470z50932 (.Y (nx2470z1), .A (nx2470z2), .B (NOT_a_1__dup_3631
           ), .C (nx52248z1)) ;
    NAND2B NOT_ix20284z49934 (.Y (nx20284z1), .A (nx20284z2), .B (nx56070z1)) ;
    NAND2B NOT_ix22498z49934 (.Y (nx22498z1), .A (nx22498z2), .B (nx32220z1)) ;
    NAND3C NOT_ix65280z50932 (.Y (nx65280z1), .A (nx6418z1), .B (
           NOT_a_1__dup_3625), .C (nx10562z1)) ;
    NAND2B NOT_ix23010z49934 (.Y (nx23010z1), .A (nx12192z1), .B (nx23010z2)) ;
    NAND3C NOT_ix19772z50932 (.Y (nx19772z1), .A (nx34946z1), .B (nx35506z3), .C (
           nx19772z2)) ;
    NAND3C NOT_ix46881z50932 (.Y (nx46881z1), .A (nx7836z1), .B (nx52784z3), .C (
           nx46881z2)) ;
    NAND3C NOT_ix60450z50932 (.Y (nx60450z1), .A (nx14918z1), .B (nx55534z2), .C (
           nx60450z2)) ;
    NAND3C NOT_ix27840z50932 (.Y (nx27840z1), .A (nx49501z1), .B (nx32756z2), .C (
           nx27840z2)) ;
    NAND3C NOT_ix14942z50932 (.Y (nx14942z1), .A (nx39776z1), .B (nx55510z2), .C (
           nx14942z2)) ;
    NAND3C NOT_ix7812z50932 (.Y (nx7812z1), .A (nx3006z1), .B (nx52808z2), .C (
           nx7812z2)) ;
    NAND3C NOT_ix34970z50932 (.Y (nx34970z1), .A (nx19748z1), .B (nx35482z2), .C (
           nx34970z2)) ;
    NAND3C NOT_ix12216z50932 (.Y (nx12216z1), .A (nx11298z1), .B (nx8409z1), .C (
           nx12216z2)) ;
    NAND3C NOT_ix10538z50932 (.Y (nx10538z1), .A (NOT_a_0__dup_3648), .B (
           nx10538z2), .C (NOT_a_1__dup_3647)) ;
    NAND3C NOT_ix32244z50932 (.Y (nx32244z1), .A (NOT_a_0__dup_3653), .B (
           nx32244z2), .C (NOT_a_1__dup_3652)) ;
    NAND3C NOT_ix56046z50932 (.Y (nx56046z1), .A (NOT_a_0__dup_3658), .B (
           nx56046z2), .C (NOT_a_1__dup_3657)) ;
    NAND3C NOT_ix8373z50932 (.Y (nx8373z1), .A (NOT_a_1__dup_3631), .B (
           NOT_a_0__dup_3632), .C (nx8373z2)) ;
    NAND3C NOT_ix15368z50932 (.Y (nx15368z1), .A (nx15368z2), .B (
           NOT_a_1__dup_3637), .C (NOT_a_0__dup_3638)) ;
    NAND3C NOT_ix27414z50932 (.Y (nx27414z1), .A (NOT_a_0_), .B (NOT_a_1_), .C (
           nx27414z2)) ;
    NAND3C NOT_ix60876z50932 (.Y (nx60876z1), .A (NOT_a_1__dup_3625), .B (
           NOT_a_0__dup_3626), .C (nx60876z2)) ;
    XA1B sclear_and_0_dup_114_rename981 (.Y (sclear_and_0_dup_114), .A (
         ENCR_DEV_encry_cnt[0]), .B (ENCR_DEV_prev[2]), .C (nx63528z1)) ;
    XA1C sclear_and_1_dup_115_rename982 (.Y (sclear_and_1_dup_115), .A (
         ENCR_DEV_encry_cnt[1]), .B (nx24762z1), .C (nx63528z1)) ;
    XA1C sclear_and_2_dup_116_rename983 (.Y (sclear_and_2_dup_116), .A (
         nx18020z1), .B (ENCR_DEV_encry_cnt[2]), .C (nx63528z1)) ;
    AND3B sclear_and_3_dup_117_rename984 (.Y (sclear_and_3_dup_117), .A (
          ENCR_DEV_prev_6__int), .B (ENCR_DEV_prev[3]), .C (inc_d_3__dup_2781)
          ) ;
    XA1C sclear_and_4_dup_118_rename985 (.Y (sclear_and_4_dup_118), .A (
         nx38048z1), .B (ENCR_DEV_encry_cnt[4]), .C (nx63528z1)) ;
    AND3B sclear_and_5_dup_119_rename986 (.Y (sclear_and_5_dup_119), .A (
          ENCR_DEV_prev_6__int), .B (ENCR_DEV_prev[3]), .C (inc_d_5__dup_2783)
          ) ;
    XA1C sclear_and_6_dup_120_rename987 (.Y (sclear_and_6_dup_120), .A (
         ENCR_DEV_encry_cnt[6]), .B (nx57089z1), .C (nx63528z1)) ;
    XA1C sclear_and_7_dup_121_rename988 (.Y (sclear_and_7_dup_121), .A (
         ENCR_DEV_encry_cnt[7]), .B (nx31201z1), .C (nx63528z1)) ;
    AND3B sclear_and_8_dup_122_rename989 (.Y (sclear_and_8_dup_122), .A (
          ENCR_DEV_prev_6__int), .B (ENCR_DEV_prev[3]), .C (inc_d_8__dup_2786)
          ) ;
    NAND2 NOT_ix52196z24339 (.Y (nx52196z2), .A (ENCR_DEV_encry_cnt[5]), .B (
          ENCR_DEV_encry_cnt[4])) ;
    NAND2 NOT_ix24762z24338 (.Y (nx24762z1), .A (ENCR_DEV_prev[2]), .B (
          ENCR_DEV_encry_cnt[0])) ;
    NAND3 NOT_ix18020z24337 (.Y (nx18020z1), .A (ENCR_DEV_prev[2]), .B (
          ENCR_DEV_encry_cnt[0]), .C (ENCR_DEV_encry_cnt[1])) ;
    NAND3A NOT_ix38048z50930 (.Y (nx38048z1), .A (nx18020z1), .B (
           ENCR_DEV_encry_cnt[3]), .C (ENCR_DEV_encry_cnt[2])) ;
    NAND3A NOT_ix52196z50930 (.Y (nx52196z1), .A (nx52196z2), .B (
           ENCR_DEV_encry_cnt[7]), .C (ENCR_DEV_encry_cnt[6])) ;
    NAND3A NOT_ix57089z50930 (.Y (nx57089z1), .A (nx38048z1), .B (
           ENCR_DEV_encry_cnt[5]), .C (ENCR_DEV_encry_cnt[4])) ;
    NAND3B NOT_ix31201z50931 (.Y (nx31201z1), .A (nx38048z1), .B (nx52196z2), .C (
           ENCR_DEV_encry_cnt[6])) ;
    AX1 inc_d_3__dup_2781_rename990 (.Y (inc_d_3__dup_2781), .A (nx18020z1), .B (
        ENCR_DEV_encry_cnt[2]), .C (ENCR_DEV_encry_cnt[3])) ;
    AX1 inc_d_5__dup_2783_rename991 (.Y (inc_d_5__dup_2783), .A (nx38048z1), .B (
        ENCR_DEV_encry_cnt[4]), .C (ENCR_DEV_encry_cnt[5])) ;
    AX1B inc_d_8__dup_2786_rename992 (.Y (inc_d_8__dup_2786), .A (nx38048z1), .B (
         nx52196z1), .C (ENCR_DEV_encry_cnt[8])) ;
    NAND3A NOT_ix32158z50930 (.Y (nx32158z1), .A (NOT_FIFO_DEV_rtlc5n43_int), .B (
           FIFO_DEV_rtlc_wadd_n4[0]), .C (FIFO_DEV_rtlc_wadd_n4[1])) ;
    AX1C inc_d_0__dup_2797_rename993 (.Y (inc_d_0__dup_2797), .A (WRITE), .B (
         NOT_CONDITION_0_), .C (FIFO_DEV_rtlc_wadd_n4[0])) ;
    AX1 inc_d_1__dup_2798_rename994 (.Y (inc_d_1__dup_2798), .A (
        NOT_FIFO_DEV_rtlc5n43_int), .B (FIFO_DEV_rtlc_wadd_n4[0]), .C (
        FIFO_DEV_rtlc_wadd_n4[1])) ;
    XNOR2 inc_d_2__dup_2799_rename995 (.Y (inc_d_2__dup_2799), .A (
          FIFO_DEV_rtlc_wadd_n4[2]), .B (nx32158z1)) ;
    AX1 inc_d_3__dup_2800_rename996 (.Y (inc_d_3__dup_2800), .A (nx32158z1), .B (
        FIFO_DEV_rtlc_wadd_n4[2]), .C (FIFO_DEV_rtlc_wadd_n4[3])) ;
    AX1B inc_d_4__dup_2801_rename997 (.Y (inc_d_4__dup_2801), .A (nx49948z1), .B (
         nx32158z1), .C (FIFO_DEV_rtlc_wadd_n4[4])) ;
    AX1B inc_d_5__dup_2802_rename998 (.Y (inc_d_5__dup_2802), .A (nx32158z1), .B (
         nx32158z3), .C (FIFO_DEV_rtlc_wadd_n4[5])) ;
    AX1B inc_d_6__dup_2803_rename999 (.Y (inc_d_6__dup_2803), .A (nx32158z1), .B (
         nx16808z1), .C (FIFO_DEV_rtlc_wadd_n4[6])) ;
    AX1B inc_d_7__dup_2804_rename1000 (.Y (inc_d_7__dup_2804), .A (nx65298z1), .B (
         nx32158z1), .C (FIFO_DEV_rtlc_wadd_n4[7])) ;
    AOI1D ix54164z47392 (.Y (nx54164z2), .A (FIFO_DEV_count[3]), .B (
          FIFO_DEV_count[2]), .C (READ_int)) ;
    AOI1D ix50324z47393 (.Y (nx50324z3), .A (FIFO_DEV_count[5]), .B (
          FIFO_DEV_count[4]), .C (READ_int)) ;
    AO1 ix57994z5368 (.Y (nx57994z3), .A (FIFO_DEV_count[6]), .B (READ_int), .C (
        nx50324z3)) ;
    MAJ3 a_0__dup_274_rename1001 (.Y (a_0__dup_274), .A (FIFO_DEV_count[1]), .B (
         FIFO_DEV_count[0]), .C (READ_int)) ;
    MAJ3 ix47598z58058 (.Y (nx47598z1), .A (FIFO_DEV_count[2]), .B (READ_int), .C (
         a_0__dup_274)) ;
    AO1A a_0__dup_276_rename1002 (.Y (a_0__dup_276), .A (nx54164z1), .B (
         a_0__dup_274), .C (nx54164z2)) ;
    MAJ3 ix27570z58058 (.Y (nx27570z1), .A (FIFO_DEV_count[4]), .B (READ_int), .C (
         a_0__dup_276)) ;
    AO1A ix50324z40555 (.Y (nx50324z1), .A (nx50324z2), .B (a_0__dup_276), .C (
         nx50324z3)) ;
    AO1A ix57994z40555 (.Y (nx57994z1), .A (nx57994z2), .B (a_0__dup_276), .C (
         nx57994z3)) ;
    AOI5 NOT_ix50324z64472 (.Y (nx50324z2), .A (READ_int), .C (FIFO_DEV_count[5]
         ), .B (FIFO_DEV_count[4])) ;
    INV a_0__dup_2819_rename1003 (.Y (a_0__dup_2819), .A (FIFO_DEV_count[0])) ;
    AOI5 NOT_ix54164z64471 (.Y (nx54164z1), .A (READ_int), .C (FIFO_DEV_count[3]
         ), .B (FIFO_DEV_count[2])) ;
    XO1A NOT_ix57994z43527 (.Y (nx57994z2), .A (FIFO_DEV_count[6]), .B (READ_int
         ), .C (nx50324z2)) ;
    XOR3 incdec_mux_1_dup_99_rename1004 (.Y (incdec_mux_1_dup_99), .A (
         FIFO_DEV_count[1]), .B (FIFO_DEV_count[0]), .C (READ_int)) ;
    XOR3 incdec_mux_2_dup_100_rename1005 (.Y (incdec_mux_2_dup_100), .A (
         FIFO_DEV_count[2]), .B (READ_int), .C (a_0__dup_274)) ;
    XOR3 incdec_mux_3_dup_101_rename1006 (.Y (incdec_mux_3_dup_101), .A (
         FIFO_DEV_count[3]), .B (READ_int), .C (nx47598z1)) ;
    XOR3 incdec_mux_4_dup_102_rename1007 (.Y (incdec_mux_4_dup_102), .A (
         FIFO_DEV_count[4]), .B (READ_int), .C (a_0__dup_276)) ;
    XOR3 incdec_mux_5_dup_103_rename1008 (.Y (incdec_mux_5_dup_103), .A (
         FIFO_DEV_count[5]), .B (READ_int), .C (nx27570z1)) ;
    XOR3 incdec_mux_6_dup_104_rename1009 (.Y (incdec_mux_6_dup_104), .A (
         FIFO_DEV_count[6]), .B (READ_int), .C (nx50324z1)) ;
    XOR3 incdec_mux_7_dup_105_rename1010 (.Y (incdec_mux_7_dup_105), .A (
         FIFO_DEV_count[7]), .B (READ_int), .C (nx57994z1)) ;
    NAND2B ENCR_DEV_rtlc15_2329_or_250_ix23410z49934 (.Y (nx23410z1), .A (
           ENCR_DEV_prev_1___repl0), .B (ENCR_DEV_prev[2])) ;
    NAND2B ENCR_DEV_rtlc15_2329_or_250_ix3438z49937 (.Y (nx3438z4), .A (
           ENCR_DEV_prev[8]), .B (ENCR_DEV_prev_6__int)) ;
    NAND3B NOT_ENCR_DEV_rtlc_835_and_296_ix10507z50932 (.Y (nx10507z2), .A (
           STB_KEY_int), .B (nx9510z3), .C (ENCR_DEV_prev[2])) ;
    NAND2A NOT_ENCR_DEV_rtlc_839_and_297_ix9510z49942 (.Y (nx9510z10), .A (
           STB_KEY_int), .B (ENCR_DEV_prev[8])) ;
    NAND3A NOT_ENCR_DEV_rtlc_841_and_298_ix9510z50931 (.Y (nx9510z2), .A (
           STB_KEY_int), .B (ENCR_DEV_prev[2]), .C (nx9510z3)) ;
    AO1C ENCR_DEV_rtlc_842_or_299_ix9510z40564 (.Y (nx9510z8), .A (CONDITION_1_)
         , .B (ENCR_DEV_prev[3]), .C (nx9510z9)) ;
    NAND2A NOT_ENCR_DEV_rtlc_851_and_300_ix36622z49934 (.Y (nx36622z2), .A (
           STB_KEY_int), .B (ENCR_DEV_prev_1___repl0)) ;
    AO1B NOT_ENCR_DEV_rtlc_863_and_302_ix3438z40557 (.Y (nx3438z2), .A (
         ENCR_DEV_prev[4]), .B (STB_DATA_int), .C (STB_KEY_int)) ;
    NAND3B NOT_ENCR_DEV_rtlc_1093_and_303_ix18636z50932 (.Y (nx18636z2), .A (
           ENCR_DEV_prev[8]), .B (ENCR_DEV_prev[3]), .C (nx45632z3)) ;
    AND2B ENCR_DEV_modgen_counter_key_cnt_ix45632z1960 (.Y (nx45632z1), .A (
          ENCR_DEV_rtlc12_X_0_n169), .B (ENCR_DEV_key_cnt[0])) ;
    XA1B ENCR_DEV_modgen_counter_key_cnt_ix44635z21033 (.Y (nx44635z1), .A (
         ENCR_DEV_key_cnt[1]), .B (ENCR_DEV_key_cnt[0]), .C (
         ENCR_DEV_rtlc12_X_0_n169)) ;
    XA1C ENCR_DEV_modgen_counter_key_cnt_ix43638z21034 (.Y (nx43638z1), .A (
         ENCR_DEV_key_cnt[2]), .B (nx43638z2), .C (ENCR_DEV_rtlc12_X_0_n169)) ;
    XA1C ENCR_DEV_modgen_counter_key_cnt_ix42641z21034 (.Y (nx42641z1), .A (
         nx40647z3), .B (ENCR_DEV_key_cnt[3]), .C (ENCR_DEV_rtlc12_X_0_n169)) ;
    XA1C ENCR_DEV_modgen_counter_key_cnt_ix41644z21034 (.Y (nx41644z1), .A (
         nx39650z3), .B (ENCR_DEV_key_cnt[4]), .C (ENCR_DEV_rtlc12_X_0_n169)) ;
    XA1C ENCR_DEV_modgen_counter_key_cnt_ix40647z21034 (.Y (nx40647z1), .A (
         nx40647z2), .B (ENCR_DEV_key_cnt[5]), .C (ENCR_DEV_rtlc12_X_0_n169)) ;
    XA1C ENCR_DEV_modgen_counter_key_cnt_ix39650z21034 (.Y (nx39650z1), .A (
         nx39650z2), .B (ENCR_DEV_key_cnt[6]), .C (ENCR_DEV_rtlc12_X_0_n169)) ;
    NAND2 NOT_ENCR_DEV_modgen_counter_key_cnt_inc_ix43638z24339 (.Y (nx43638z2)
          , .A (ENCR_DEV_key_cnt[1]), .B (ENCR_DEV_key_cnt[0])) ;
    NAND3 NOT_ENCR_DEV_modgen_counter_key_cnt_inc_ix40647z24339 (.Y (nx40647z3)
          , .A (ENCR_DEV_key_cnt[2]), .B (ENCR_DEV_key_cnt[1]), .C (
          ENCR_DEV_key_cnt[0])) ;
    NAND3A NOT_ENCR_DEV_modgen_counter_key_cnt_inc_ix39650z50932 (.Y (nx39650z3)
           , .A (nx43638z2), .B (ENCR_DEV_key_cnt[2]), .C (ENCR_DEV_key_cnt[3])
           ) ;
    NAND3A NOT_ENCR_DEV_modgen_counter_key_cnt_inc_ix40647z50931 (.Y (nx40647z2)
           , .A (nx40647z3), .B (ENCR_DEV_key_cnt[3]), .C (ENCR_DEV_key_cnt[4])
           ) ;
    NAND3A NOT_ENCR_DEV_modgen_counter_key_cnt_inc_ix39650z50931 (.Y (nx39650z2)
           , .A (nx39650z3), .B (ENCR_DEV_key_cnt[4]), .C (ENCR_DEV_key_cnt[5])
           ) ;
    NAND3C ENCR_DEV_modgen_or_0_ix15492z50935 (.Y (nx15492z4), .A (
           ENCR_DEV_cnt_init[8]), .B (ENCR_DEV_cnt_init[7]), .C (
           ENCR_DEV_cnt_init[9])) ;
    MX2C FIFO_DEV_rtlc14_20_or_596_ix59980z26291 (.Y (nx59980z1), .A (
         NOT_CONDITION_0_), .S (READ_int), .B (CONDITION_1_)) ;
    NAND3A FIFO_DEV_ix0_cmp_240__ix37353z50931 (.Y (nx37353z2), .A (nx37353z3), 
           .B (FIFO_DEV_rtlc_wadd_n4[7]), .C (FIFO_DEV_rtlc_wadd_n4[6])) ;
    NAND3B FIFO_DEV_ix0_cmp_224__ix19403z50932 (.Y (nx19403z2), .A (nx19403z3), 
           .B (FIFO_DEV_rtlc_wadd_n4[4]), .C (FIFO_DEV_rtlc_wadd_n4[5])) ;
    NAND3B FIFO_DEV_ix0_cmp_208__ix2452z50932 (.Y (nx2452z2), .A (nx19403z3), .B (
           FIFO_DEV_rtlc_wadd_n4[5]), .C (FIFO_DEV_rtlc_wadd_n4[4])) ;
    NAND2 FIFO_DEV_ix0_cmp_192__ix19403z24340 (.Y (nx19403z3), .A (
          FIFO_DEV_rtlc_wadd_n4[7]), .B (FIFO_DEV_rtlc_wadd_n4[6])) ;
    NAND3C FIFO_DEV_ix0_cmp_192__ix50038z50933 (.Y (nx50038z2), .A (nx19403z3), 
           .B (FIFO_DEV_rtlc_wadd_n4[5]), .C (FIFO_DEV_rtlc_wadd_n4[4])) ;
    NAND3B FIFO_DEV_ix0_cmp_176__ix45412z50932 (.Y (nx45412z2), .A (
           FIFO_DEV_rtlc_wadd_n4[6]), .B (nx37353z3), .C (
           FIFO_DEV_rtlc_wadd_n4[7])) ;
    NAND3B FIFO_DEV_ix0_cmp_160__ix63362z50932 (.Y (nx63362z2), .A (
           FIFO_DEV_rtlc_wadd_n4[4]), .B (nx63362z3), .C (
           FIFO_DEV_rtlc_wadd_n4[5])) ;
    NAND3B FIFO_DEV_ix0_cmp_144__ix15776z50932 (.Y (nx15776z2), .A (
           FIFO_DEV_rtlc_wadd_n4[5]), .B (nx63362z3), .C (
           FIFO_DEV_rtlc_wadd_n4[4])) ;
    NAND2A FIFO_DEV_ix0_cmp_128__ix63362z49935 (.Y (nx63362z3), .A (
           FIFO_DEV_rtlc_wadd_n4[6]), .B (FIFO_DEV_rtlc_wadd_n4[7])) ;
    NAND3C FIFO_DEV_ix0_cmp_128__ix32727z50933 (.Y (nx32727z2), .A (
           FIFO_DEV_rtlc_wadd_n4[5]), .B (FIFO_DEV_rtlc_wadd_n4[4]), .C (
           nx63362z3)) ;
    NAND3B FIFO_DEV_ix0_cmp_112__ix50677z50932 (.Y (nx50677z2), .A (
           FIFO_DEV_rtlc_wadd_n4[7]), .B (nx37353z3), .C (
           FIFO_DEV_rtlc_wadd_n4[6])) ;
    NAND3B FIFO_DEV_ix0_cmp_96__ix2092z50932 (.Y (nx2092z2), .A (nx2092z3), .B (
           FIFO_DEV_rtlc_wadd_n4[4]), .C (FIFO_DEV_rtlc_wadd_n4[5])) ;
    NAND3B FIFO_DEV_ix0_cmp_80__ix9565z50932 (.Y (nx9565z2), .A (nx2092z3), .B (
           FIFO_DEV_rtlc_wadd_n4[5]), .C (FIFO_DEV_rtlc_wadd_n4[4])) ;
    NAND2A FIFO_DEV_ix0_cmp_64__ix2092z49935 (.Y (nx2092z3), .A (
           FIFO_DEV_rtlc_wadd_n4[7]), .B (FIFO_DEV_rtlc_wadd_n4[6])) ;
    NAND3C FIFO_DEV_ix0_cmp_64__ix27515z50933 (.Y (nx27515z2), .A (nx2092z3), .B (
           FIFO_DEV_rtlc_wadd_n4[5]), .C (FIFO_DEV_rtlc_wadd_n4[4])) ;
    NAND2 FIFO_DEV_ix0_cmp_48__ix37353z24340 (.Y (nx37353z3), .A (
          FIFO_DEV_rtlc_wadd_n4[5]), .B (FIFO_DEV_rtlc_wadd_n4[4])) ;
    NAND3C FIFO_DEV_ix0_cmp_48__ix44466z50933 (.Y (nx44466z2), .A (
           FIFO_DEV_rtlc_wadd_n4[7]), .B (FIFO_DEV_rtlc_wadd_n4[6]), .C (
           nx37353z3)) ;
    NAND2A FIFO_DEV_ix0_cmp_32__ix62416z49935 (.Y (nx62416z3), .A (
           FIFO_DEV_rtlc_wadd_n4[4]), .B (FIFO_DEV_rtlc_wadd_n4[5])) ;
    NAND3C FIFO_DEV_ix0_cmp_32__ix62416z50933 (.Y (nx62416z2), .A (
           FIFO_DEV_rtlc_wadd_n4[7]), .B (FIFO_DEV_rtlc_wadd_n4[6]), .C (
           nx62416z3)) ;
    NAND2A FIFO_DEV_ix0_cmp_16__ix13831z49935 (.Y (nx13831z3), .A (
           FIFO_DEV_rtlc_wadd_n4[5]), .B (FIFO_DEV_rtlc_wadd_n4[4])) ;
    NAND3C FIFO_DEV_ix0_cmp_16__ix13831z50933 (.Y (nx13831z2), .A (
           FIFO_DEV_rtlc_wadd_n4[7]), .B (FIFO_DEV_rtlc_wadd_n4[6]), .C (
           nx13831z3)) ;
    NAND3A FIFO_DEV_ix0_cmp_15__ix37353z50933 (.Y (nx37353z4), .A (nx49948z1), .B (
           FIFO_DEV_rtlc_wadd_n4[1]), .C (FIFO_DEV_rtlc_wadd_n4[0])) ;
    NAND3B FIFO_DEV_ix0_cmp_14__ix36356z50932 (.Y (nx36356z2), .A (nx49948z1), .B (
           FIFO_DEV_rtlc_wadd_n4[0]), .C (FIFO_DEV_rtlc_wadd_n4[1])) ;
    NAND3B FIFO_DEV_ix0_cmp_13__ix35359z50932 (.Y (nx35359z2), .A (nx49948z1), .B (
           FIFO_DEV_rtlc_wadd_n4[1]), .C (FIFO_DEV_rtlc_wadd_n4[0])) ;
    NAND2 FIFO_DEV_ix0_cmp_12__ix49948z24338 (.Y (nx49948z1), .A (
          FIFO_DEV_rtlc_wadd_n4[3]), .B (FIFO_DEV_rtlc_wadd_n4[2])) ;
    NAND3C FIFO_DEV_ix0_cmp_12__ix34362z50933 (.Y (nx34362z2), .A (nx49948z1), .B (
           FIFO_DEV_rtlc_wadd_n4[1]), .C (FIFO_DEV_rtlc_wadd_n4[0])) ;
    NAND3B FIFO_DEV_ix0_cmp_11__ix33365z50932 (.Y (nx33365z2), .A (
           FIFO_DEV_rtlc_wadd_n4[2]), .B (nx33365z3), .C (
           FIFO_DEV_rtlc_wadd_n4[3])) ;
    NAND3B FIFO_DEV_ix0_cmp_10__ix32368z50932 (.Y (nx32368z2), .A (
           FIFO_DEV_rtlc_wadd_n4[0]), .B (nx32368z3), .C (
           FIFO_DEV_rtlc_wadd_n4[1])) ;
    NAND3B FIFO_DEV_ix0_cmp_9__ix30372z50932 (.Y (nx30372z2), .A (
           FIFO_DEV_rtlc_wadd_n4[1]), .B (nx32368z3), .C (
           FIFO_DEV_rtlc_wadd_n4[0])) ;
    NAND2A FIFO_DEV_ix0_cmp_8__ix32368z49935 (.Y (nx32368z3), .A (
           FIFO_DEV_rtlc_wadd_n4[2]), .B (FIFO_DEV_rtlc_wadd_n4[3])) ;
    NAND3C FIFO_DEV_ix0_cmp_8__ix29375z50933 (.Y (nx29375z2), .A (
           FIFO_DEV_rtlc_wadd_n4[1]), .B (FIFO_DEV_rtlc_wadd_n4[0]), .C (
           nx32368z3)) ;
    NAND3B FIFO_DEV_ix0_cmp_7__ix28378z50932 (.Y (nx28378z2), .A (
           FIFO_DEV_rtlc_wadd_n4[3]), .B (nx33365z3), .C (
           FIFO_DEV_rtlc_wadd_n4[2])) ;
    NAND3B FIFO_DEV_ix0_cmp_6__ix27381z50932 (.Y (nx27381z2), .A (
           FIFO_DEV_rtlc_wadd_n4[0]), .B (nx27381z3), .C (
           FIFO_DEV_rtlc_wadd_n4[1])) ;
    NAND3B FIFO_DEV_ix0_cmp_5__ix26384z50932 (.Y (nx26384z2), .A (
           FIFO_DEV_rtlc_wadd_n4[1]), .B (nx27381z3), .C (
           FIFO_DEV_rtlc_wadd_n4[0])) ;
    NAND2A FIFO_DEV_ix0_cmp_4__ix27381z49935 (.Y (nx27381z3), .A (
           FIFO_DEV_rtlc_wadd_n4[3]), .B (FIFO_DEV_rtlc_wadd_n4[2])) ;
    NAND3C FIFO_DEV_ix0_cmp_4__ix25387z50933 (.Y (nx25387z2), .A (
           FIFO_DEV_rtlc_wadd_n4[1]), .B (FIFO_DEV_rtlc_wadd_n4[0]), .C (
           nx27381z3)) ;
    NAND2 FIFO_DEV_ix0_cmp_3__ix33365z24340 (.Y (nx33365z3), .A (
          FIFO_DEV_rtlc_wadd_n4[1]), .B (FIFO_DEV_rtlc_wadd_n4[0])) ;
    NAND3C FIFO_DEV_ix0_cmp_3__ix24390z50933 (.Y (nx24390z2), .A (
           FIFO_DEV_rtlc_wadd_n4[3]), .B (FIFO_DEV_rtlc_wadd_n4[2]), .C (
           nx33365z3)) ;
    NAND2A FIFO_DEV_ix0_cmp_2__ix23393z49935 (.Y (nx23393z3), .A (
           FIFO_DEV_rtlc_wadd_n4[0]), .B (FIFO_DEV_rtlc_wadd_n4[1])) ;
    NAND3C FIFO_DEV_ix0_cmp_2__ix23393z50933 (.Y (nx23393z2), .A (
           FIFO_DEV_rtlc_wadd_n4[3]), .B (FIFO_DEV_rtlc_wadd_n4[2]), .C (
           nx23393z3)) ;
    NAND2A FIFO_DEV_ix0_cmp_1__ix22396z49935 (.Y (nx22396z3), .A (
           FIFO_DEV_rtlc_wadd_n4[1]), .B (FIFO_DEV_rtlc_wadd_n4[0])) ;
    NAND3C FIFO_DEV_ix0_cmp_1__ix22396z50933 (.Y (nx22396z2), .A (
           FIFO_DEV_rtlc_wadd_n4[3]), .B (FIFO_DEV_rtlc_wadd_n4[2]), .C (
           nx22396z3)) ;
    NAND2B FIFO_DEV_ix0_cmp_0__ix21399z49936 (.Y (nx21399z3), .A (
           FIFO_DEV_rtlc_wadd_n4[1]), .B (FIFO_DEV_rtlc_wadd_n4[0])) ;
    NAND3C FIFO_DEV_ix0_cmp_0__ix21399z50933 (.Y (nx21399z2), .A (
           FIFO_DEV_rtlc_wadd_n4[3]), .B (FIFO_DEV_rtlc_wadd_n4[2]), .C (
           nx21399z3)) ;
    NAND2B FIFO_DEV_ix0_cmp_0__ix31781z49936 (.Y (nx31781z3), .A (
           FIFO_DEV_rtlc_wadd_n4[5]), .B (FIFO_DEV_rtlc_wadd_n4[4])) ;
    NAND3C FIFO_DEV_ix0_cmp_0__ix31781z50933 (.Y (nx31781z2), .A (
           FIFO_DEV_rtlc_wadd_n4[7]), .B (FIFO_DEV_rtlc_wadd_n4[6]), .C (
           nx31781z3)) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_0__ix35840z14896 (.Y (
        nx35840z1), .A (ENCR_DEV_t_3[7]), .S (b_0__int), .B (ENCR_DEV_t_3[0])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_1__ix36837z14896 (.Y (
        nx36837z1), .A (ENCR_DEV_t_3[6]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[0])) ;
    NAND2A NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_1__ix36837z49934
            (.Y (nx36837z2), .A (b_0__int), .B (ENCR_DEV_key_reg[3])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_2__ix37834z14896 (.Y (
        nx37834z1), .A (ENCR_DEV_t_3[5]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[1])) ;
    NAND2A NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_2__ix37834z49934
            (.Y (nx37834z2), .A (b_0__int), .B (ENCR_DEV_key_reg[4])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_3__ix38831z14896 (.Y (
        nx38831z1), .A (ENCR_DEV_t_3[4]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[2])) ;
    NAND2A NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_3__ix38831z49934
            (.Y (nx38831z2), .A (b_0__int), .B (ENCR_DEV_key_reg[5])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_4__ix39828z14896 (.Y (
        nx39828z1), .A (ENCR_DEV_t_3[3]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[3])) ;
    NAND2A NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_4__ix39828z49934
            (.Y (nx39828z2), .A (b_0__int), .B (ENCR_DEV_key_reg[6])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_5__ix40825z14896 (.Y (
        nx40825z1), .A (ENCR_DEV_t_3[2]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[4])) ;
    NAND2A NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_5__ix40825z49934
            (.Y (nx40825z2), .A (b_0__int), .B (ENCR_DEV_key_reg[7])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_6__ix41822z14896 (.Y (
        nx41822z1), .A (ENCR_DEV_t_3[1]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[5])) ;
    NAND2A NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_6__ix41822z49934
            (.Y (nx41822z2), .A (b_0__int), .B (ENCR_DEV_key_reg[8])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_7__ix42819z14896 (.Y (
        nx42819z1), .A (ENCR_DEV_t_3[0]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[6])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_8__ix43816z14896 (.Y (
        nx43816z1), .A (ENCR_DEV_reg_str_1[0]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[7])) ;
    NAND2A NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_8__ix43816z49934
            (.Y (nx43816z2), .A (b_0__int), .B (ENCR_DEV_key_reg[10])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_9__ix44813z14896 (.Y (
        nx44813z1), .A (ENCR_DEV_reg_str_1[1]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[8])) ;
    NAND2A NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_9__ix44813z49934
            (.Y (nx44813z2), .A (b_0__int), .B (ENCR_DEV_key_reg[11])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_10__ix32187z14896 (.Y (
        nx32187z1), .A (ENCR_DEV_reg_str_1[2]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[9])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_10__ix32187z49934
            (.Y (nx32187z2), .A (b_0__int), .B (ENCR_DEV_key_reg[12])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_11__ix31190z14896 (.Y (
        nx31190z1), .A (ENCR_DEV_reg_str_1[3]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[10])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_11__ix31190z49934
            (.Y (nx31190z2), .A (b_0__int), .B (ENCR_DEV_key_reg[13])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_12__ix30193z14896 (.Y (
        nx30193z1), .A (ENCR_DEV_reg_str_1[4]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[11])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_12__ix30193z49934
            (.Y (nx30193z2), .A (b_0__int), .B (ENCR_DEV_key_reg[14])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_13__ix29196z14896 (.Y (
        nx29196z1), .A (ENCR_DEV_reg_str_1[5]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[12])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_13__ix29196z49934
            (.Y (nx29196z2), .A (b_0__int), .B (ENCR_DEV_key_reg[15])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_14__ix28199z14896 (.Y (
        nx28199z1), .A (ENCR_DEV_reg_str_1[6]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[13])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_14__ix28199z49934
            (.Y (nx28199z2), .A (b_0__int), .B (ENCR_DEV_key_reg[16])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_15__ix27202z14896 (.Y (
        nx27202z1), .A (ENCR_DEV_reg_str_1[7]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[14])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_15__ix27202z49934
            (.Y (nx27202z2), .A (b_0__int), .B (ENCR_DEV_key_reg[17])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_16__ix26205z14896 (.Y (
        nx26205z1), .A (ENCR_DEV_reg_str_1[8]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[15])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_16__ix26205z49934
            (.Y (nx26205z2), .A (b_0__int), .B (ENCR_DEV_key_reg[18])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_17__ix25208z14896 (.Y (
        nx25208z1), .A (ENCR_DEV_reg_str_1[9]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[16])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_17__ix25208z49934
            (.Y (nx25208z2), .A (b_0__int), .B (ENCR_DEV_key_reg[19])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_18__ix24211z14896 (.Y (
        nx24211z1), .A (ENCR_DEV_reg_str_1[10]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[17])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_18__ix24211z49934
            (.Y (nx24211z2), .A (b_0__int), .B (ENCR_DEV_key_reg[20])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_19__ix23214z14896 (.Y (
        nx23214z1), .A (ENCR_DEV_reg_str_1[11]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[18])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_19__ix23214z49934
            (.Y (nx23214z2), .A (b_0__int), .B (ENCR_DEV_key_reg[21])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_20__ix21218z14896 (.Y (
        nx21218z1), .A (ENCR_DEV_reg_str_1[12]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[19])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_20__ix21218z49934
            (.Y (nx21218z2), .A (b_0__int), .B (ENCR_DEV_key_reg[22])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_21__ix20221z14896 (.Y (
        nx20221z1), .A (ENCR_DEV_reg_str_1[13]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[20])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_21__ix20221z49934
            (.Y (nx20221z2), .A (b_0__int), .B (ENCR_DEV_key_reg[23])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_22__ix19224z14896 (.Y (
        nx19224z1), .A (ENCR_DEV_reg_str_1[14]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[21])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_22__ix19224z49934
            (.Y (nx19224z2), .A (b_0__int), .B (ENCR_DEV_key_reg[24])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_23__ix18227z14896 (.Y (
        nx18227z1), .A (ENCR_DEV_reg_str_1[15]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[22])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_23__ix18227z49934
            (.Y (nx18227z2), .A (b_0__int), .B (ENCR_DEV_key_reg[25])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_24__ix17230z14896 (.Y (
        nx17230z1), .A (ENCR_DEV_reg_str_1[16]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[23])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_24__ix17230z49934
            (.Y (nx17230z2), .A (b_0__int), .B (ENCR_DEV_key_reg[26])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_25__ix16233z14896 (.Y (
        nx16233z1), .A (ENCR_DEV_reg_str_1[17]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[24])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_25__ix16233z49934
            (.Y (nx16233z2), .A (b_0__int), .B (ENCR_DEV_key_reg[27])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_26__ix15236z14896 (.Y (
        nx15236z1), .A (ENCR_DEV_reg_str_1[18]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[25])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_26__ix15236z49934
            (.Y (nx15236z2), .A (b_0__int), .B (ENCR_DEV_key_reg[28])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_27__ix14239z14896 (.Y (
        nx14239z1), .A (ENCR_DEV_reg_str_1[19]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[26])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_27__ix14239z49934
            (.Y (nx14239z2), .A (b_0__int), .B (ENCR_DEV_key_reg[29])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_28__ix13242z14896 (.Y (
        nx13242z1), .A (ENCR_DEV_reg_str_1[20]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[27])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_28__ix13242z49934
            (.Y (nx13242z2), .A (b_0__int), .B (ENCR_DEV_key_reg[30])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_29__ix12245z14896 (.Y (
        nx12245z1), .A (ENCR_DEV_reg_str_1[21]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[28])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_29__ix12245z49934
            (.Y (nx12245z2), .A (b_0__int), .B (ENCR_DEV_key_reg[31])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_30__ix10249z14896 (.Y (
        nx10249z1), .A (ENCR_DEV_reg_str_1[22]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[29])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_30__ix10249z49934
            (.Y (nx10249z2), .A (b_0__int), .B (ENCR_DEV_key_reg[32])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_31__ix9252z14896 (.Y (
        nx9252z1), .A (ENCR_DEV_reg_str_1[23]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[30])) ;
    NAND2A NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_31__ix9252z49934
            (.Y (nx9252z2), .A (b_0__int), .B (ENCR_DEV_key_reg[33])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_32__ix8255z14896 (.Y (
        nx8255z1), .A (ENCR_DEV_reg_str_1[24]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[31])) ;
    NAND2A NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_32__ix8255z49934
            (.Y (nx8255z2), .A (b_0__int), .B (ENCR_DEV_key_reg[34])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_33__ix7258z14896 (.Y (
        nx7258z1), .A (ENCR_DEV_reg_str_1[25]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[32])) ;
    NAND2A NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_33__ix7258z49934
            (.Y (nx7258z2), .A (b_0__int), .B (ENCR_DEV_key_reg[35])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_34__ix6261z14896 (.Y (
        nx6261z1), .A (ENCR_DEV_reg_str_1[26]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[33])) ;
    NAND2A NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_34__ix6261z49934
            (.Y (nx6261z2), .A (b_0__int), .B (ENCR_DEV_key_reg[36])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_35__ix5264z14896 (.Y (
        nx5264z1), .A (ENCR_DEV_reg_str_1[27]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[34])) ;
    NAND2A NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_35__ix5264z49934
            (.Y (nx5264z2), .A (b_0__int), .B (ENCR_DEV_key_reg[37])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_36__ix4267z14896 (.Y (
        nx4267z1), .A (ENCR_DEV_reg_str_1[28]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[35])) ;
    NAND2A NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_36__ix4267z49934
            (.Y (nx4267z2), .A (b_0__int), .B (ENCR_DEV_key_reg[38])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_37__ix3270z14896 (.Y (
        nx3270z1), .A (ENCR_DEV_reg_str_1[29]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[36])) ;
    NAND2A NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_37__ix3270z49934
            (.Y (nx3270z2), .A (b_0__int), .B (ENCR_DEV_key_reg[39])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_38__ix2273z14896 (.Y (
        nx2273z1), .A (ENCR_DEV_reg_str_1[30]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[37])) ;
    NAND2A NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_38__ix2273z49934
            (.Y (nx2273z2), .A (b_0__int), .B (ENCR_DEV_key_reg[40])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_39__ix1276z14896 (.Y (
        nx1276z1), .A (ENCR_DEV_reg_str_1[31]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[38])) ;
    NAND2A NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_39__ix1276z49934
            (.Y (nx1276z2), .A (b_0__int), .B (ENCR_DEV_key_reg[41])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_40__ix64816z14896 (.Y (
        nx64816z1), .A (ENCR_DEV_reg_str_1[32]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[39])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_40__ix64816z49934
            (.Y (nx64816z2), .A (b_0__int), .B (ENCR_DEV_key_reg[42])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_41__ix63819z14896 (.Y (
        nx63819z1), .A (ENCR_DEV_reg_str_1[33]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[40])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_41__ix63819z49934
            (.Y (nx63819z2), .A (b_0__int), .B (ENCR_DEV_key_reg[43])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_42__ix62822z14896 (.Y (
        nx62822z1), .A (ENCR_DEV_reg_str_1[34]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[41])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_42__ix62822z49934
            (.Y (nx62822z2), .A (b_0__int), .B (ENCR_DEV_key_reg[44])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_43__ix61825z14896 (.Y (
        nx61825z1), .A (ENCR_DEV_reg_str_1[35]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[42])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_43__ix61825z49934
            (.Y (nx61825z2), .A (b_0__int), .B (ENCR_DEV_key_reg[45])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_44__ix60828z14896 (.Y (
        nx60828z1), .A (ENCR_DEV_reg_str_1[36]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[43])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_44__ix60828z49934
            (.Y (nx60828z2), .A (b_0__int), .B (ENCR_DEV_key_reg[46])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_45__ix59831z14896 (.Y (
        nx59831z1), .A (ENCR_DEV_reg_str_1[37]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[44])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_45__ix59831z49934
            (.Y (nx59831z2), .A (b_0__int), .B (ENCR_DEV_key_reg[47])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_46__ix58834z14896 (.Y (
        nx58834z1), .A (ENCR_DEV_reg_str_1[38]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[45])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_46__ix58834z49934
            (.Y (nx58834z2), .A (b_0__int), .B (ENCR_DEV_key_reg[48])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_47__ix57837z14896 (.Y (
        nx57837z1), .A (ENCR_DEV_reg_str_1[39]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[46])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_47__ix57837z49934
            (.Y (nx57837z2), .A (b_0__int), .B (ENCR_DEV_key_reg[49])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_48__ix56840z14896 (.Y (
        nx56840z1), .A (ENCR_DEV_reg_str_1[40]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[47])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_48__ix56840z49934
            (.Y (nx56840z2), .A (b_0__int), .B (ENCR_DEV_key_reg[50])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_49__ix55843z14896 (.Y (
        nx55843z1), .A (ENCR_DEV_reg_str_1[41]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[48])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_49__ix55843z49934
            (.Y (nx55843z2), .A (b_0__int), .B (ENCR_DEV_key_reg[51])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_50__ix53847z14896 (.Y (
        nx53847z1), .A (ENCR_DEV_reg_str_1[42]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[49])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_50__ix53847z49934
            (.Y (nx53847z2), .A (b_0__int), .B (ENCR_DEV_key_reg[52])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_51__ix52850z14896 (.Y (
        nx52850z1), .A (ENCR_DEV_reg_str_1[43]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[50])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_51__ix52850z49934
            (.Y (nx52850z2), .A (b_0__int), .B (ENCR_DEV_key_reg[53])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_52__ix51853z14896 (.Y (
        nx51853z1), .A (ENCR_DEV_reg_str_1[44]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[51])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_52__ix51853z49934
            (.Y (nx51853z2), .A (b_0__int), .B (ENCR_DEV_key_reg[54])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_53__ix50856z14896 (.Y (
        nx50856z1), .A (ENCR_DEV_reg_str_1[45]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[52])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_53__ix50856z49934
            (.Y (nx50856z2), .A (b_0__int), .B (ENCR_DEV_key_reg[55])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_54__ix49859z14896 (.Y (
        nx49859z1), .A (ENCR_DEV_reg_str_1[46]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[53])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_54__ix49859z49934
            (.Y (nx49859z2), .A (b_0__int), .B (ENCR_DEV_key_reg[56])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_55__ix48862z14896 (.Y (
        nx48862z1), .A (ENCR_DEV_reg_str_1[47]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[54])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_55__ix48862z49934
            (.Y (nx48862z2), .A (b_0__int), .B (ENCR_DEV_key_reg[57])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_56__ix47865z14896 (.Y (
        nx47865z1), .A (ENCR_DEV_reg_str_1[48]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[55])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_56__ix47865z49934
            (.Y (nx47865z2), .A (b_0__int), .B (ENCR_DEV_key_reg[58])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_57__ix46868z14896 (.Y (
        nx46868z1), .A (ENCR_DEV_reg_str_1[49]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[56])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_57__ix46868z49934
            (.Y (nx46868z2), .A (b_0__int), .B (ENCR_DEV_key_reg[59])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_58__ix45871z14896 (.Y (
        nx45871z1), .A (ENCR_DEV_reg_str_1[50]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[57])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_58__ix45871z49934
            (.Y (nx45871z2), .A (b_0__int), .B (ENCR_DEV_key_reg[60])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_59__ix44874z14896 (.Y (
        nx44874z1), .A (ENCR_DEV_reg_str_1[51]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[58])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_59__ix44874z49934
            (.Y (nx44874z2), .A (b_0__int), .B (ENCR_DEV_key_reg[61])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_60__ix42878z14896 (.Y (
        nx42878z1), .A (ENCR_DEV_reg_str_1[52]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[59])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_60__ix42878z49934
            (.Y (nx42878z2), .A (b_0__int), .B (ENCR_DEV_key_reg[62])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_61__ix41881z14896 (.Y (
        nx41881z1), .A (ENCR_DEV_reg_str_1[53]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[60])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_61__ix41881z49934
            (.Y (nx41881z2), .A (b_0__int), .B (ENCR_DEV_key_reg[63])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_62__ix40884z14896 (.Y (
        nx40884z1), .A (ENCR_DEV_reg_str_1[54]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[61])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_62__ix40884z49934
            (.Y (nx40884z2), .A (b_0__int), .B (ENCR_DEV_key_reg[64])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_63__ix39887z14896 (.Y (
        nx39887z1), .A (ENCR_DEV_reg_str_1[55]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[62])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_63__ix39887z49934
            (.Y (nx39887z2), .A (b_0__int), .B (ENCR_DEV_key_reg[65])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_64__ix38890z14896 (.Y (
        nx38890z1), .A (ENCR_DEV_reg_str_1[56]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[63])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_64__ix38890z49934
            (.Y (nx38890z2), .A (b_0__int), .B (ENCR_DEV_key_reg[66])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_65__ix37893z14896 (.Y (
        nx37893z1), .A (ENCR_DEV_reg_str_1[57]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[64])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_65__ix37893z49934
            (.Y (nx37893z2), .A (b_0__int), .B (ENCR_DEV_key_reg[67])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_66__ix36896z14896 (.Y (
        nx36896z1), .A (ENCR_DEV_reg_str_1[58]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[65])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_66__ix36896z49934
            (.Y (nx36896z2), .A (b_0__int), .B (ENCR_DEV_key_reg[68])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_67__ix35899z14896 (.Y (
        nx35899z1), .A (ENCR_DEV_reg_str_1[59]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[66])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_67__ix35899z49934
            (.Y (nx35899z2), .A (b_0__int), .B (ENCR_DEV_key_reg[69])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_68__ix34902z14896 (.Y (
        nx34902z1), .A (ENCR_DEV_reg_str_1[60]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[67])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_68__ix34902z49934
            (.Y (nx34902z2), .A (b_0__int), .B (ENCR_DEV_key_reg[70])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_69__ix33905z14896 (.Y (
        nx33905z1), .A (ENCR_DEV_reg_str_1[61]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[68])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_69__ix33905z49934
            (.Y (nx33905z2), .A (b_0__int), .B (ENCR_DEV_key_reg[71])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_70__ix31909z14896 (.Y (
        nx31909z1), .A (ENCR_DEV_reg_str_1[62]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[69])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_70__ix31909z49934
            (.Y (nx31909z2), .A (b_0__int), .B (ENCR_DEV_key_reg[72])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_71__ix30912z14896 (.Y (
        nx30912z1), .A (ENCR_DEV_reg_str_1[63]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[70])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_71__ix30912z49934
            (.Y (nx30912z2), .A (b_0__int), .B (ENCR_DEV_key_reg[73])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_72__ix29915z14896 (.Y (
        nx29915z1), .A (ENCR_DEV_reg_str_1[64]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[71])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_72__ix29915z49934
            (.Y (nx29915z2), .A (b_0__int), .B (ENCR_DEV_key_reg[74])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_73__ix28918z14896 (.Y (
        nx28918z1), .A (ENCR_DEV_reg_str_1[65]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[72])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_73__ix28918z49934
            (.Y (nx28918z2), .A (b_0__int), .B (ENCR_DEV_key_reg[75])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_74__ix27921z14896 (.Y (
        nx27921z1), .A (ENCR_DEV_reg_str_1[66]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[73])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_74__ix27921z49934
            (.Y (nx27921z2), .A (b_0__int), .B (ENCR_DEV_key_reg[76])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_75__ix26924z14896 (.Y (
        nx26924z1), .A (ENCR_DEV_reg_str_1[67]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[74])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_75__ix26924z49934
            (.Y (nx26924z2), .A (b_0__int), .B (ENCR_DEV_key_reg[77])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_76__ix25927z14896 (.Y (
        nx25927z1), .A (ENCR_DEV_reg_str_1[68]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[75])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_76__ix25927z49934
            (.Y (nx25927z2), .A (b_0__int), .B (ENCR_DEV_key_reg[78])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_77__ix24930z14896 (.Y (
        nx24930z1), .A (ENCR_DEV_reg_str_1[69]), .S (b_0__int), .B (
        ENCR_DEV_reg_str_1[76])) ;
    NAND2A 
           NOT_prec_sel2mux_ENCR_DEV_reg_str_1_select_15i1Bus15_77__ix24930z49934
            (.Y (nx24930z2), .A (b_0__int), .B (ENCR_DEV_key_reg[79])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i79Bus16_78__ix23933z14896 (.Y (
        nx23933z1), .A (ENCR_DEV_reg_str_1[70]), .S (ENCR_DEV_prev[8]), .B (
        ENCR_DEV_reg_str_1[77])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i79Bus16_79__ix22936z14896 (.Y (
        nx22936z1), .A (ENCR_DEV_reg_str_1[71]), .S (ENCR_DEV_prev[8]), .B (
        ENCR_DEV_reg_str_1[78])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i79Bus16_80__ix20940z14896 (.Y (
        nx20940z1), .A (ENCR_DEV_reg_str_1[72]), .S (ENCR_DEV_prev[8]), .B (
        ENCR_DEV_reg_str_1[79])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i79Bus16_81__ix19943z14896 (.Y (
        nx19943z1), .A (ENCR_DEV_reg_str_1[73]), .S (ENCR_DEV_prev[8]), .B (
        ENCR_DEV_reg_str_1[80])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i79Bus16_82__ix18946z14896 (.Y (
        nx18946z1), .A (ENCR_DEV_reg_str_1[74]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_1[81])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i79Bus16_83__ix17949z14896 (.Y (
        nx17949z1), .A (ENCR_DEV_reg_str_1[75]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_1[82])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i79Bus16_84__ix16952z14896 (.Y (
        nx16952z1), .A (ENCR_DEV_reg_str_1[76]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_1[83])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i79Bus16_85__ix15955z14896 (.Y (
        nx15955z1), .A (ENCR_DEV_reg_str_1[77]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_1[84])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i79Bus16_86__ix14958z14896 (.Y (
        nx14958z1), .A (ENCR_DEV_reg_str_1[78]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_1[85])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i79Bus16_87__ix13961z14896 (.Y (
        nx13961z1), .A (ENCR_DEV_reg_str_1[79]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_1[86])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i79Bus16_88__ix12964z14896 (.Y (
        nx12964z1), .A (ENCR_DEV_reg_str_1[80]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_1[87])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i79Bus16_89__ix11967z14896 (.Y (
        nx11967z1), .A (ENCR_DEV_reg_str_1[81]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_1[88])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i79Bus16_90__ix9971z14896 (.Y (
        nx9971z1), .A (ENCR_DEV_reg_str_1[82]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_1[89])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i79Bus16_91__ix8974z14896 (.Y (
        nx8974z1), .A (ENCR_DEV_reg_str_1[83]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_1[90])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_1_select_15i79Bus16_92__ix7977z14896 (.Y (
        nx7977z1), .A (ENCR_DEV_reg_str_1[84]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_1[91])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i130Bus39_80__ix58629z14896 (.Y (
        nx58629z1), .A (ENCR_DEV_reg_str_2[72]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_2[79])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i130Bus39_81__ix59626z14896 (.Y (
        nx59626z1), .A (ENCR_DEV_reg_str_2[73]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_2[80])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i130Bus39_82__ix60623z14896 (.Y (
        nx60623z1), .A (ENCR_DEV_reg_str_2[74]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_2[81])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i130Bus39_83__ix61620z14896 (.Y (
        nx61620z1), .A (ENCR_DEV_reg_str_2[75]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_2[82])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_0__ix21254z14896 (.Y (
        nx21254z1), .A (ENCR_DEV_t_2[7]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_t_2[0])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_1__ix20257z14896 (.Y (
        nx20257z1), .A (ENCR_DEV_t_2[6]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_3[0])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_2__ix19260z14896 (.Y (
        nx19260z1), .A (ENCR_DEV_t_2[5]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_3[1])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_3__ix18263z14896 (.Y (
        nx18263z1), .A (ENCR_DEV_t_2[4]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_3[2])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_4__ix17266z14896 (.Y (
        nx17266z1), .A (ENCR_DEV_t_2[3]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_3[3])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_5__ix16269z14896 (.Y (
        nx16269z1), .A (ENCR_DEV_t_2[2]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_3[4])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_6__ix15272z14896 (.Y (
        nx15272z1), .A (ENCR_DEV_t_2[1]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_3[5])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_7__ix14275z14896 (.Y (
        nx14275z1), .A (ENCR_DEV_t_2[0]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_3[6])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_8__ix13278z14896 (.Y (
        nx13278z1), .A (ENCR_DEV_reg_str_3[0]), .S (ENCR_DEV_prev_8___repl6), .B (
        ENCR_DEV_reg_str_3[7])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_9__ix12281z14896 (.Y (
        nx12281z1), .A (ENCR_DEV_reg_str_3[1]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[8])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_10__ix4121z14896 (.Y (
        nx4121z1), .A (ENCR_DEV_reg_str_3[2]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[9])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_11__ix3124z14896 (.Y (
        nx3124z1), .A (ENCR_DEV_reg_str_3[3]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[10])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_12__ix2127z14896 (.Y (
        nx2127z1), .A (ENCR_DEV_reg_str_3[4]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[11])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_13__ix1130z14896 (.Y (
        nx1130z1), .A (ENCR_DEV_reg_str_3[5]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[12])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_14__ix133z14896 (.Y (
        nx133z1), .A (ENCR_DEV_reg_str_3[6]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[13])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_15__ix64672z14896 (.Y (
        nx64672z1), .A (ENCR_DEV_reg_str_3[7]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[14])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_16__ix63675z14896 (.Y (
        nx63675z1), .A (ENCR_DEV_reg_str_3[8]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[15])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_17__ix62678z14896 (.Y (
        nx62678z1), .A (ENCR_DEV_reg_str_3[9]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[16])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_18__ix61681z14896 (.Y (
        nx61681z1), .A (ENCR_DEV_reg_str_3[10]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[17])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_19__ix60684z14896 (.Y (
        nx60684z1), .A (ENCR_DEV_reg_str_3[11]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[18])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_20__ix58688z14896 (.Y (
        nx58688z1), .A (ENCR_DEV_reg_str_3[12]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[19])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_21__ix57691z14896 (.Y (
        nx57691z1), .A (ENCR_DEV_reg_str_3[13]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[20])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_22__ix56694z14896 (.Y (
        nx56694z1), .A (ENCR_DEV_reg_str_3[14]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[21])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_23__ix55697z14896 (.Y (
        nx55697z1), .A (ENCR_DEV_reg_str_3[15]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[22])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_24__ix54700z14896 (.Y (
        nx54700z1), .A (ENCR_DEV_reg_str_3[16]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[23])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_25__ix53703z14896 (.Y (
        nx53703z1), .A (ENCR_DEV_reg_str_3[17]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[24])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_26__ix52706z14896 (.Y (
        nx52706z1), .A (ENCR_DEV_reg_str_3[18]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[25])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_27__ix51709z14896 (.Y (
        nx51709z1), .A (ENCR_DEV_reg_str_3[19]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[26])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_28__ix50712z14896 (.Y (
        nx50712z1), .A (ENCR_DEV_reg_str_3[20]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[27])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_29__ix49715z14896 (.Y (
        nx49715z1), .A (ENCR_DEV_reg_str_3[21]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[28])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_30__ix47719z14896 (.Y (
        nx47719z1), .A (ENCR_DEV_reg_str_3[22]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[29])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_31__ix46722z14896 (.Y (
        nx46722z1), .A (ENCR_DEV_reg_str_3[23]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[30])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_32__ix45725z14896 (.Y (
        nx45725z1), .A (ENCR_DEV_reg_str_3[24]), .S (ENCR_DEV_prev_8___repl5), .B (
        ENCR_DEV_reg_str_3[31])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_33__ix44728z14896 (.Y (
        nx44728z1), .A (ENCR_DEV_reg_str_3[25]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[32])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_34__ix43731z14896 (.Y (
        nx43731z1), .A (ENCR_DEV_reg_str_3[26]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[33])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_35__ix42734z14896 (.Y (
        nx42734z1), .A (ENCR_DEV_reg_str_3[27]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[34])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_36__ix41737z14896 (.Y (
        nx41737z1), .A (ENCR_DEV_reg_str_3[28]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[35])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_37__ix40740z14896 (.Y (
        nx40740z1), .A (ENCR_DEV_reg_str_3[29]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[36])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_38__ix39743z14896 (.Y (
        nx39743z1), .A (ENCR_DEV_reg_str_3[30]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[37])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_39__ix38746z14896 (.Y (
        nx38746z1), .A (ENCR_DEV_reg_str_3[31]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[38])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_40__ix36750z14896 (.Y (
        nx36750z1), .A (ENCR_DEV_reg_str_3[32]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[39])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_41__ix35753z14896 (.Y (
        nx35753z1), .A (ENCR_DEV_reg_str_3[33]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[40])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_42__ix34756z14896 (.Y (
        nx34756z1), .A (ENCR_DEV_reg_str_3[34]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[41])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_43__ix33759z14896 (.Y (
        nx33759z1), .A (ENCR_DEV_reg_str_3[35]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[42])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_44__ix32762z14896 (.Y (
        nx32762z1), .A (ENCR_DEV_reg_str_3[36]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[43])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_45__ix31765z14896 (.Y (
        nx31765z1), .A (ENCR_DEV_reg_str_3[37]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[44])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_46__ix30768z14896 (.Y (
        nx30768z1), .A (ENCR_DEV_reg_str_3[38]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[45])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_47__ix29771z14896 (.Y (
        nx29771z1), .A (ENCR_DEV_reg_str_3[39]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[46])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_48__ix28774z14896 (.Y (
        nx28774z1), .A (ENCR_DEV_reg_str_3[40]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[47])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_49__ix27777z14896 (.Y (
        nx27777z1), .A (ENCR_DEV_reg_str_3[41]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[48])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_50__ix25781z14896 (.Y (
        nx25781z1), .A (ENCR_DEV_reg_str_3[42]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[49])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_51__ix24784z14896 (.Y (
        nx24784z1), .A (ENCR_DEV_reg_str_3[43]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[50])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_52__ix23787z14896 (.Y (
        nx23787z1), .A (ENCR_DEV_reg_str_3[44]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[51])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_53__ix22790z14896 (.Y (
        nx22790z1), .A (ENCR_DEV_reg_str_3[45]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[52])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_54__ix21793z14896 (.Y (
        nx21793z1), .A (ENCR_DEV_reg_str_3[46]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[53])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_55__ix20796z14896 (.Y (
        nx20796z1), .A (ENCR_DEV_reg_str_3[47]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[54])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_56__ix19799z14896 (.Y (
        nx19799z1), .A (ENCR_DEV_reg_str_3[48]), .S (ENCR_DEV_prev_8___repl4), .B (
        ENCR_DEV_reg_str_3[55])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_57__ix18802z14896 (.Y (
        nx18802z1), .A (ENCR_DEV_reg_str_3[49]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[56])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_58__ix17805z14896 (.Y (
        nx17805z1), .A (ENCR_DEV_reg_str_3[50]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[57])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_59__ix16808z14896 (.Y (
        nx16808z2), .A (ENCR_DEV_reg_str_3[51]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[58])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_60__ix14812z14896 (.Y (
        nx14812z1), .A (ENCR_DEV_reg_str_3[52]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[59])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_61__ix13815z14896 (.Y (
        nx13815z1), .A (ENCR_DEV_reg_str_3[53]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[60])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_62__ix12818z14896 (.Y (
        nx12818z1), .A (ENCR_DEV_reg_str_3[54]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[61])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_63__ix11821z14896 (.Y (
        nx11821z1), .A (ENCR_DEV_reg_str_3[55]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[62])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_64__ix10824z14896 (.Y (
        nx10824z1), .A (ENCR_DEV_reg_str_3[56]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[63])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_65__ix9827z14896 (.Y (
        nx9827z1), .A (ENCR_DEV_reg_str_3[57]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[64])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_66__ix8830z14896 (.Y (
        nx8830z1), .A (ENCR_DEV_reg_str_3[58]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[65])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_67__ix7833z14896 (.Y (
        nx7833z1), .A (ENCR_DEV_reg_str_3[59]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[66])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_68__ix6836z14896 (.Y (
        nx6836z1), .A (ENCR_DEV_reg_str_3[60]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[67])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_69__ix5839z14896 (.Y (
        nx5839z1), .A (ENCR_DEV_reg_str_3[61]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[68])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_70__ix3843z14896 (.Y (
        nx3843z1), .A (ENCR_DEV_reg_str_3[62]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[69])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_71__ix2846z14896 (.Y (
        nx2846z1), .A (ENCR_DEV_reg_str_3[63]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[70])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_72__ix1849z14896 (.Y (
        nx1849z1), .A (ENCR_DEV_reg_str_3[64]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[71])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_73__ix852z14896 (.Y (
        nx852z1), .A (ENCR_DEV_reg_str_3[65]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[72])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_74__ix65391z14896 (.Y (
        nx65391z1), .A (ENCR_DEV_reg_str_3[66]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[73])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_75__ix64394z14896 (.Y (
        nx64394z1), .A (ENCR_DEV_reg_str_3[67]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[74])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_76__ix63397z14896 (.Y (
        nx63397z1), .A (ENCR_DEV_reg_str_3[68]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[75])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_77__ix62400z14896 (.Y (
        nx62400z1), .A (ENCR_DEV_reg_str_3[69]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[76])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_78__ix61403z14896 (.Y (
        nx61403z1), .A (ENCR_DEV_reg_str_3[70]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[77])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_79__ix60406z14896 (.Y (
        nx60406z1), .A (ENCR_DEV_reg_str_3[71]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[78])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_80__ix58410z14896 (.Y (
        nx58410z1), .A (ENCR_DEV_reg_str_3[72]), .S (ENCR_DEV_prev_8___repl3), .B (
        ENCR_DEV_reg_str_3[79])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_81__ix57413z14896 (.Y (
        nx57413z1), .A (ENCR_DEV_reg_str_3[73]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[80])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_82__ix56416z14896 (.Y (
        nx56416z1), .A (ENCR_DEV_reg_str_3[74]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[81])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_83__ix55419z14896 (.Y (
        nx55419z1), .A (ENCR_DEV_reg_str_3[75]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[82])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_84__ix54422z14896 (.Y (
        nx54422z1), .A (ENCR_DEV_reg_str_3[76]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[83])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_85__ix53425z14896 (.Y (
        nx53425z1), .A (ENCR_DEV_reg_str_3[77]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[84])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_86__ix52428z14896 (.Y (
        nx52428z1), .A (ENCR_DEV_reg_str_3[78]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[85])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_87__ix51431z14896 (.Y (
        nx51431z1), .A (ENCR_DEV_reg_str_3[79]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[86])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_88__ix50434z14896 (.Y (
        nx50434z1), .A (ENCR_DEV_reg_str_3[80]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[87])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_89__ix49437z14896 (.Y (
        nx49437z1), .A (ENCR_DEV_reg_str_3[81]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[88])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_90__ix47441z14896 (.Y (
        nx47441z1), .A (ENCR_DEV_reg_str_3[82]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[89])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_91__ix46444z14896 (.Y (
        nx46444z1), .A (ENCR_DEV_reg_str_3[83]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[90])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_92__ix45447z14896 (.Y (
        nx45447z1), .A (ENCR_DEV_reg_str_3[84]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[91])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_93__ix44450z14896 (.Y (
        nx44450z1), .A (ENCR_DEV_reg_str_3[85]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[92])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_94__ix43453z14896 (.Y (
        nx43453z1), .A (ENCR_DEV_reg_str_3[86]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[93])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_95__ix42456z14896 (.Y (
        nx42456z1), .A (ENCR_DEV_reg_str_3[87]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[94])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_96__ix41459z14896 (.Y (
        nx41459z1), .A (ENCR_DEV_reg_str_3[88]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[95])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_97__ix40462z14896 (.Y (
        nx40462z1), .A (ENCR_DEV_reg_str_3[89]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[96])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_98__ix39465z14896 (.Y (
        nx39465z1), .A (ENCR_DEV_reg_str_3[90]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[97])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_99__ix38468z14896 (.Y (
        nx38468z1), .A (ENCR_DEV_reg_str_3[91]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[98])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_100__ix27151z14896 (.Y (
        nx27151z1), .A (ENCR_DEV_reg_str_3[92]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[99])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_101__ix28148z14896 (.Y (
        nx28148z1), .A (ENCR_DEV_reg_str_3[93]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[100])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_102__ix29145z14896 (.Y (
        nx29145z1), .A (ENCR_DEV_reg_str_3[94]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[101])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_103__ix30142z14896 (.Y (
        nx30142z1), .A (ENCR_DEV_reg_str_3[95]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[102])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_104__ix31139z14896 (.Y (
        nx31139z1), .A (ENCR_DEV_reg_str_3[96]), .S (ENCR_DEV_prev_8___repl2), .B (
        ENCR_DEV_reg_str_3[103])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_105__ix32136z14896 (.Y (
        nx32136z1), .A (ENCR_DEV_reg_str_3[97]), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_3[104])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_106__ix33133z14896 (.Y (
        nx33133z1), .A (ENCR_DEV_reg_str_3[98]), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_3[105])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_3_select_15i134Bus40_107__ix34130z14896 (.Y (
        nx34130z1), .A (ENCR_DEV_reg_str_3[99]), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_3[106])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i245Bus17_1__ix24478z14896 (.Y (
        nx24478z1), .A (ENCR_DEV_t_1_6_), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[0])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i245Bus17_2__ix23481z14896 (.Y (
        nx23481z1), .A (ENCR_DEV_t_1_5_), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[1])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i247Bus18_4__ix21487z14896 (.Y (
        nx21487z1), .A (ENCR_DEV_t_1_3_), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[3])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i247Bus18_5__ix20490z14896 (.Y (
        nx20490z1), .A (ENCR_DEV_t_1_2_), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[4])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i247Bus18_6__ix19493z14896 (.Y (
        nx19493z1), .A (ENCR_DEV_t_1_1_), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[5])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i247Bus18_7__ix18496z14896 (.Y (
        nx18496z1), .A (ENCR_DEV_t_1_0_), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[6])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i251_ix16502z14896 (.Y (
        nx16502z1), .A (ENCR_DEV_reg_str_2[1]), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[8])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i252Bus19_11__ix48379z14896 (.Y (
        nx48379z1), .A (ENCR_DEV_reg_str_2[3]), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[10])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i252Bus19_12__ix49376z14896 (.Y (
        nx49376z1), .A (ENCR_DEV_reg_str_2[4]), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[11])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i254Bus21_15__ix52367z14896 (.Y (
        nx52367z1), .A (ENCR_DEV_reg_str_2[7]), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[14])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i254Bus21_16__ix53364z14896 (.Y (
        nx53364z1), .A (ENCR_DEV_reg_str_2[8]), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[15])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i256Bus23_19__ix56355z14896 (.Y (
        nx56355z1), .A (ENCR_DEV_reg_str_2[11]), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[18])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i256Bus23_20__ix58351z14896 (.Y (
        nx58351z1), .A (ENCR_DEV_reg_str_2[12]), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[19])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i256Bus23_21__ix59348z14896 (.Y (
        nx59348z1), .A (ENCR_DEV_reg_str_2[13]), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[20])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i259Bus24_23__ix61342z14896 (.Y (
        nx61342z1), .A (ENCR_DEV_reg_str_2[15]), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[22])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i259Bus24_24__ix62339z14896 (.Y (
        nx62339z1), .A (ENCR_DEV_reg_str_2[16]), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[23])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i259Bus24_25__ix63336z14896 (.Y (
        nx63336z1), .A (ENCR_DEV_reg_str_2[17]), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[24])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i259Bus24_26__ix64333z14896 (.Y (
        nx64333z1), .A (ENCR_DEV_reg_str_2[18]), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[25])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i259Bus24_27__ix65330z14896 (.Y (
        nx65330z1), .A (ENCR_DEV_reg_str_2[19]), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[26])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i264Bus26_31__ix4781z14896 (.Y (
        nx4781z1), .A (ENCR_DEV_reg_str_2[23]), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[30])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i264Bus26_32__ix5778z14896 (.Y (
        nx5778z1), .A (ENCR_DEV_reg_str_2[24]), .S (ENCR_DEV_prev_8___repl1), .B (
        ENCR_DEV_reg_str_2[31])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i264Bus26_33__ix6775z14896 (.Y (
        nx6775z1), .A (ENCR_DEV_reg_str_2[25]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[32])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i267_ix8769z14896 (.Y (nx8769z1
        ), .A (ENCR_DEV_reg_str_2[27]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[34])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i268_ix10763z14896 (.Y (
        nx10763z1), .A (ENCR_DEV_reg_str_2[29]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[36])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i269_ix14753z14896 (.Y (
        nx14753z1), .A (ENCR_DEV_reg_str_2[32]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[39])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i270_ix17744z14896 (.Y (
        nx17744z1), .A (ENCR_DEV_reg_str_2[35]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[42])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i271_ix19738z14896 (.Y (
        nx19738z1), .A (ENCR_DEV_reg_str_2[37]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[44])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i272_ix21732z14896 (.Y (
        nx21732z1), .A (ENCR_DEV_reg_str_2[39]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[46])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i273_ix25722z14896 (.Y (
        nx25722z1), .A (ENCR_DEV_reg_str_2[42]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[49])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i274_ix28713z14896 (.Y (
        nx28713z1), .A (ENCR_DEV_reg_str_2[45]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[52])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i275_ix30707z14896 (.Y (
        nx30707z1), .A (ENCR_DEV_reg_str_2[47]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[54])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i276Bus31_57__ix32701z14896 (.Y (
        nx32701z1), .A (ENCR_DEV_reg_str_2[49]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[56])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i276Bus31_58__ix33698z14896 (.Y (
        nx33698z1), .A (ENCR_DEV_reg_str_2[50]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[57])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i276Bus31_59__ix34695z14896 (.Y (
        nx34695z1), .A (ENCR_DEV_reg_str_2[51]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[58])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i279Bus33_63__ix39682z14896 (.Y (
        nx39682z1), .A (ENCR_DEV_reg_str_2[55]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[62])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i279Bus33_64__ix40679z14896 (.Y (
        nx40679z1), .A (ENCR_DEV_reg_str_2[56]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[63])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i281Bus35_67__ix43670z14896 (.Y (
        nx43670z1), .A (ENCR_DEV_reg_str_2[59]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[66])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i281Bus35_68__ix44667z14896 (.Y (
        nx44667z1), .A (ENCR_DEV_reg_str_2[60]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[67])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i281Bus35_69__ix45664z14896 (.Y (
        nx45664z1), .A (ENCR_DEV_reg_str_2[61]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[68])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i281Bus35_70__ix47660z14896 (.Y (
        nx47660z1), .A (ENCR_DEV_reg_str_2[62]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[69])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i285_ix49654z14896 (.Y (
        nx49654z1), .A (ENCR_DEV_reg_str_2[64]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[71])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i286Bus37_75__ix52645z14896 (.Y (
        nx52645z1), .A (ENCR_DEV_reg_str_2[67]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[74])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i286Bus37_76__ix53642z14896 (.Y (
        nx53642z1), .A (ENCR_DEV_reg_str_2[68]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[75])) ;
    MX2 prec_sel2mux_ENCR_DEV_reg_str_2_select_15i286Bus37_77__ix54639z14896 (.Y (
        nx54639z1), .A (ENCR_DEV_reg_str_2[69]), .S (ENCR_DEV_prev_8___repl0), .B (
        ENCR_DEV_reg_str_2[76])) ;
    NAND3A NOT_a_2__dup_4701_rename1011 (.Y (NOT_a_2__dup_4701), .A (
           NOT_a_4__dup_3628), .B (ENCR_DEV_err_cnt[59]), .C (
           ENCR_DEV_err_cnt[58])) ;
    NAND2B NOT_a_1__dup_4702_rename1012 (.Y (NOT_a_1__dup_4702), .A (
           NOT_a_3__dup_3640), .B (NOT_a_3__dup_3629)) ;
    NAND3C NOT_modgen_and_324_ix12216z50933 (.Y (nx12216z2), .A (
           NOT_a_1__dup_3642), .B (NOT_a_2__dup_3641), .C (NOT_a_1__dup_4702)) ;
    NAND2 NOT_modgen_and_380_ix15492z24343 (.Y (nx15492z6), .A (
          ENCR_DEV_cnt_init[4]), .B (ENCR_DEV_cnt_init[2])) ;
    NAND2 NOT_modgen_and_380_ix15492z24344 (.Y (nx15492z7), .A (
          ENCR_DEV_cnt_init[5]), .B (ENCR_DEV_cnt_init[1])) ;
    NAND3 NOT_modgen_and_380_ix15492z24354 (.Y (nx15492z8), .A (
          ENCR_DEV_cnt_init[3]), .B (ENCR_DEV_cnt_init[0]), .C (
          ENCR_DEV_cnt_init[6])) ;
    NAND2 NOT_modgen_and_381_ix9510z24342 (.Y (nx9510z5), .A (
          ENCR_DEV_encry_cnt[2]), .B (ENCR_DEV_encry_cnt[1])) ;
    NAND3A NOT_modgen_and_381_ix9510z50933 (.Y (nx9510z4), .A (nx9510z5), .B (
           ENCR_DEV_encry_cnt[4]), .C (ENCR_DEV_encry_cnt[3])) ;
    NAND2 NOT_modgen_and_381_ix9510z24344 (.Y (nx9510z7), .A (
          ENCR_DEV_encry_cnt[6]), .B (ENCR_DEV_encry_cnt[5])) ;
    NAND3B NOT_modgen_and_381_ix9510z50936 (.Y (nx9510z6), .A (nx9510z7), .B (
           ENCR_DEV_encry_cnt[8]), .C (ENCR_DEV_encry_cnt[7])) ;
    NAND3 NOT_modgen_and_382_ix11504z24346 (.Y (nx11504z9), .A (
          ENCR_DEV_err_cnt[3]), .B (ENCR_DEV_err_cnt[2]), .C (
          ENCR_DEV_err_cnt[1])) ;
    NAND3C NOT_modgen_and_382_ix11504z50940 (.Y (nx11504z8), .A (nx11298z2), .B (
           nx11298z3), .C (nx11504z9)) ;
    NAND3C NOT_modgen_and_382_ix10507z50935 (.Y (nx10507z4), .A (nx8409z2), .B (
           nx11504z3), .C (nx11504z8)) ;
    NAND2 NOT_modgen_and_382_ix11504z24355 (.Y (nx11504z17), .A (
          ENCR_DEV_err_cnt[60]), .B (ENCR_DEV_err_cnt[0])) ;
    NAND3C NOT_modgen_and_382_ix11504z50948 (.Y (nx11504z16), .A (nx49501z3), .B (
           nx49501z6), .C (nx11504z17)) ;
    NAND3C NOT_modgen_and_382_ix11504z50942 (.Y (nx11504z10), .A (nx11504z11), .B (
           NOT_a_2__dup_3641), .C (nx11504z16)) ;
    NAND3C NOT_modgen_and_382_ix11504z50933 (.Y (nx11504z2), .A (NOT_a_7_), .B (
           nx11504z8), .C (nx11504z10)) ;
    NAND2 NOT_modgen_and_382_ix11504z24358 (.Y (nx11504z20), .A (
          ENCR_DEV_err_cnt[63]), .B (ENCR_DEV_err_cnt[61])) ;
    NAND2A NOT_modgen_and_382_ix11504z49954 (.Y (nx11504z21), .A (
           NOT_a_2__dup_4701), .B (ENCR_DEV_err_cnt[62])) ;
    NAND3C NOT_modgen_and_382_ix11504z50951 (.Y (nx11504z19), .A (
           NOT_a_1__dup_4702), .B (nx11504z20), .C (nx11504z21)) ;
    NAND2 NOT_modgen_and_383_ix41852z24339 (.Y (nx41852z2), .A (
          FIFO_DEV_count[1]), .B (FIFO_DEV_count[0])) ;
    NAND3A NOT_modgen_and_383_ix41852z50930 (.Y (nx41852z1), .A (nx41852z2), .B (
           FIFO_DEV_count[3]), .C (FIFO_DEV_count[2])) ;
    NAND2 NOT_modgen_and_383_ix41852z24340 (.Y (nx41852z3), .A (
          FIFO_DEV_count[5]), .B (FIFO_DEV_count[4])) ;
    NAND2 NOT_modgen_and_383_ix41852z24341 (.Y (nx41852z4), .A (
          FIFO_DEV_count[7]), .B (FIFO_DEV_count[6])) ;
    NAND2B modgen_or_384_ix54297z49935 (.Y (nx54297z2), .A (FIFO_DEV_count[7]), 
           .B (FIFO_DEV_count[6])) ;
    NAND3C modgen_or_384_ix54297z50932 (.Y (nx54297z1), .A (FIFO_DEV_count[5]), 
           .B (FIFO_DEV_count[4]), .C (nx54297z2)) ;
    NAND2B modgen_or_384_ix54297z49936 (.Y (nx54297z3), .A (FIFO_DEV_count[3]), 
           .B (FIFO_DEV_count[2])) ;
    NAND2B modgen_or_384_ix54297z49937 (.Y (nx54297z4), .A (FIFO_DEV_count[1]), 
           .B (FIFO_DEV_count[0])) ;
    XOR3 modgen_xor_385_ix48026z10877 (.Y (nx48026z1), .A (nx48026z2), .B (
         ENCR_DEV_reg_str_2[68]), .C (ENCR_DEV_data_reg[0])) ;
    XOR3 modgen_xor_385_ix48026z10879 (.Y (nx48026z3), .A (
         ENCR_DEV_reg_str_3[65]), .B (ENCR_DEV_reg_str_1[65]), .C (
         ENCR_DEV_reg_str_2[83])) ;
    XOR3 modgen_xor_386_ix47029z10877 (.Y (nx47029z1), .A (nx47029z2), .B (
         ENCR_DEV_reg_str_1[64]), .C (ENCR_DEV_data_reg[1])) ;
    XOR3 modgen_xor_386_ix47029z10879 (.Y (nx47029z3), .A (
         ENCR_DEV_reg_str_3[109]), .B (ENCR_DEV_reg_str_1[91]), .C (
         ENCR_DEV_reg_str_2[82])) ;
    XOR3 modgen_xor_387_ix46032z10877 (.Y (nx46032z1), .A (
         ENCR_DEV_reg_str_1[63]), .B (nx46032z2), .C (ENCR_DEV_data_reg[2])) ;
    XOR3 modgen_xor_387_ix46032z10879 (.Y (nx46032z3), .A (
         ENCR_DEV_reg_str_3[108]), .B (ENCR_DEV_reg_str_1[90]), .C (
         ENCR_DEV_reg_str_2[81])) ;
    XOR3 modgen_xor_388_ix45035z10877 (.Y (nx45035z1), .A (
         ENCR_DEV_reg_str_1[62]), .B (nx45035z2), .C (ENCR_DEV_data_reg[3])) ;
    XOR3 modgen_xor_388_ix45035z10879 (.Y (nx45035z3), .A (
         ENCR_DEV_reg_str_1[89]), .B (ENCR_DEV_reg_str_2[80]), .C (
         ENCR_DEV_reg_str_3[107])) ;
    XOR3 modgen_xor_389_ix44038z10877 (.Y (nx44038z1), .A (
         ENCR_DEV_reg_str_1[61]), .B (nx44038z2), .C (ENCR_DEV_data_reg[4])) ;
    XOR3 modgen_xor_389_ix44038z10879 (.Y (nx44038z3), .A (
         ENCR_DEV_reg_str_1[88]), .B (ENCR_DEV_reg_str_2[79]), .C (
         ENCR_DEV_reg_str_3[106])) ;
    XOR3 modgen_xor_390_ix43041z10877 (.Y (nx43041z1), .A (nx43041z2), .B (
         ENCR_DEV_reg_str_1[60]), .C (ENCR_DEV_data_reg[5])) ;
    XOR3 modgen_xor_390_ix43041z10879 (.Y (nx43041z3), .A (
         ENCR_DEV_reg_str_3[105]), .B (ENCR_DEV_reg_str_1[87]), .C (
         ENCR_DEV_reg_str_2[78])) ;
    XOR3 modgen_xor_391_ix42044z10877 (.Y (nx42044z1), .A (nx42044z2), .B (
         ENCR_DEV_reg_str_1[59]), .C (ENCR_DEV_data_reg[6])) ;
    XOR3 modgen_xor_391_ix42044z10879 (.Y (nx42044z3), .A (
         ENCR_DEV_reg_str_3[59]), .B (ENCR_DEV_reg_str_1[86]), .C (
         ENCR_DEV_reg_str_2[77])) ;
    XOR3 modgen_xor_392_ix41047z10877 (.Y (nx41047z1), .A (nx41047z2), .B (
         ENCR_DEV_reg_str_1[58]), .C (ENCR_DEV_data_reg[7])) ;
    XOR3 modgen_xor_392_ix41047z10879 (.Y (nx41047z3), .A (
         ENCR_DEV_reg_str_3[103]), .B (ENCR_DEV_reg_str_1[85]), .C (
         ENCR_DEV_reg_str_2[76])) ;
    NAND3B NOT_modgen_and_393_ix27414z50933 (.Y (nx27414z3), .A (NOT_a_4_), .B (
           NOT_a_3_), .C (ENCR_DEV_err_cnt[60])) ;
    NAND3B NOT_modgen_and_393_ix27414z50932 (.Y (nx27414z2), .A (NOT_a_2_), .B (
           nx27414z3), .C (ENCR_DEV_err_cnt[61])) ;
    NAND3B NOT_modgen_and_394_ix60876z50933 (.Y (nx60876z3), .A (
           NOT_a_4__dup_3622), .B (NOT_a_3__dup_3623), .C (ENCR_DEV_err_cnt[61])
           ) ;
    NAND3B NOT_modgen_and_394_ix60876z50932 (.Y (nx60876z2), .A (
           NOT_a_2__dup_3624), .B (nx60876z3), .C (ENCR_DEV_err_cnt[62])) ;
    NAND3C NOT_modgen_and_395_ix8373z50933 (.Y (nx8373z2), .A (NOT_a_2__dup_3630
           ), .B (NOT_a_3__dup_3629), .C (NOT_a_2__dup_4701)) ;
    NAND3C NOT_modgen_and_396_ix15368z50933 (.Y (nx15368z2), .A (nx15368z3), .B (
           NOT_a_3__dup_3635), .C (NOT_a_2__dup_3636)) ;
    NAND3A NOT_modgen_and_396_ix15368z50932 (.Y (nx15368z3), .A (
           NOT_a_4__dup_3622), .B (ENCR_DEV_err_cnt[58]), .C (
           ENCR_DEV_err_cnt[57])) ;
    NAND3C NOT_modgen_and_397_ix10538z50933 (.Y (nx10538z2), .A (
           NOT_a_3__dup_3635), .B (NOT_a_3__dup_3645), .C (NOT_a_2__dup_3646)) ;
    NAND3C NOT_modgen_and_398_ix32244z50933 (.Y (nx32244z2), .A (
           NOT_a_3__dup_3650), .B (NOT_a_3_), .C (NOT_a_2__dup_3651)) ;
    NAND3C NOT_modgen_and_399_ix56046z50933 (.Y (nx56046z2), .A (
           NOT_a_2__dup_3656), .B (NOT_a_3__dup_3655), .C (NOT_a_3__dup_3623)) ;
    AO1A NOT_ENCR_DEV_ix7969z40555 (.Y (nx7969z1), .A (STB_KEY_int), .B (
         nx18636z1), .C (nx18636z2)) ;
    NAND3C NOT_ENCR_DEV_ix19668z50932 (.Y (nx19668z1), .A (
           ENCR_DEV_rtlc15_PS14_n166), .B (ENCR_DEV_prev[3]), .C (
           ENCR_DEV_rtlcn483__repl0)) ;
    AO1D NOT_ENCR_DEV_ix55223z40558 (.Y (nx55223z1), .A (nx23410z1), .B (
         nx3438z4), .C (ENCR_DEV_rtlcn483__repl0)) ;
    NAND3C ENCR_DEV_rtlc15_PS14_n166_rename1013 (.Y (ENCR_DEV_rtlc15_PS14_n166)
           , .A (ENCR_DEV_prev_5___repl0), .B (ENCR_DEV_prev[4]), .C (
           ENCR_DEV_prev[0])) ;
    NAND3C NOT_FIFO_DEV_ix37353z50932 (.Y (nx37353z1), .A (nx37353z2), .B (
           nx37353z4), .C (NOT_FIFO_DEV_rtlc5n43_int)) ;
    NAND3C NOT_FIFO_DEV_ix36356z50932 (.Y (nx36356z1), .A (nx37353z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx36356z2)) ;
    NAND3C NOT_FIFO_DEV_ix35359z50932 (.Y (nx35359z1), .A (nx37353z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx35359z2)) ;
    NAND3C NOT_FIFO_DEV_ix34362z50932 (.Y (nx34362z1), .A (nx37353z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx34362z2)) ;
    NAND3C NOT_FIFO_DEV_ix33365z50932 (.Y (nx33365z1), .A (nx37353z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx33365z2)) ;
    NAND3C NOT_FIFO_DEV_ix32368z50932 (.Y (nx32368z1), .A (nx37353z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx32368z2)) ;
    NAND3C NOT_FIFO_DEV_ix30372z50932 (.Y (nx30372z1), .A (nx37353z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx30372z2)) ;
    NAND3C NOT_FIFO_DEV_ix29375z50932 (.Y (nx29375z1), .A (nx37353z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx29375z2)) ;
    NAND3C NOT_FIFO_DEV_ix28378z50932 (.Y (nx28378z1), .A (nx37353z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx28378z2)) ;
    NAND3C NOT_FIFO_DEV_ix27381z50932 (.Y (nx27381z1), .A (nx37353z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx27381z2)) ;
    NAND3C NOT_FIFO_DEV_ix26384z50932 (.Y (nx26384z1), .A (nx37353z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx26384z2)) ;
    NAND3C NOT_FIFO_DEV_ix25387z50932 (.Y (nx25387z1), .A (nx37353z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx25387z2)) ;
    NAND3C NOT_FIFO_DEV_ix24390z50932 (.Y (nx24390z1), .A (nx37353z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx24390z2)) ;
    NAND3C NOT_FIFO_DEV_ix23393z50932 (.Y (nx23393z1), .A (nx37353z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx23393z2)) ;
    NAND3C NOT_FIFO_DEV_ix22396z50932 (.Y (nx22396z1), .A (nx37353z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx22396z2)) ;
    NAND3C NOT_FIFO_DEV_ix21399z50932 (.Y (nx21399z1), .A (nx37353z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx21399z2)) ;
    NAND3C NOT_FIFO_DEV_ix19403z50932 (.Y (nx19403z1), .A (nx37353z4), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx19403z2)) ;
    NAND3C NOT_FIFO_DEV_ix18406z50932 (.Y (nx18406z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx36356z2), .C (nx19403z2)) ;
    NAND3C NOT_FIFO_DEV_ix17409z50932 (.Y (nx17409z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx35359z2), .C (nx19403z2)) ;
    NAND3C NOT_FIFO_DEV_ix16412z50932 (.Y (nx16412z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx34362z2), .C (nx19403z2)) ;
    NAND3C NOT_FIFO_DEV_ix15415z50932 (.Y (nx15415z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx33365z2), .C (nx19403z2)) ;
    NAND3C NOT_FIFO_DEV_ix14418z50932 (.Y (nx14418z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx32368z2), .C (nx19403z2)) ;
    NAND3C NOT_FIFO_DEV_ix13421z50932 (.Y (nx13421z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx30372z2), .C (nx19403z2)) ;
    NAND3C NOT_FIFO_DEV_ix12424z50932 (.Y (nx12424z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx29375z2), .C (nx19403z2)) ;
    NAND3C NOT_FIFO_DEV_ix11427z50932 (.Y (nx11427z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx28378z2), .C (nx19403z2)) ;
    NAND3C NOT_FIFO_DEV_ix10430z50932 (.Y (nx10430z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx27381z2), .C (nx19403z2)) ;
    NAND3C NOT_FIFO_DEV_ix8434z50932 (.Y (nx8434z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx26384z2), .C (nx19403z2)) ;
    NAND3C NOT_FIFO_DEV_ix7437z50932 (.Y (nx7437z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx25387z2), .C (nx19403z2)) ;
    NAND3C NOT_FIFO_DEV_ix6440z50932 (.Y (nx6440z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx24390z2), .C (nx19403z2)) ;
    NAND3C NOT_FIFO_DEV_ix5443z50932 (.Y (nx5443z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx23393z2), .C (nx19403z2)) ;
    NAND3C NOT_FIFO_DEV_ix4446z50932 (.Y (nx4446z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx22396z2), .C (nx19403z2)) ;
    NAND3C NOT_FIFO_DEV_ix3449z50932 (.Y (nx3449z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx21399z2), .C (nx19403z2)) ;
    NAND3C NOT_FIFO_DEV_ix2452z50932 (.Y (nx2452z1), .A (nx37353z4), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx2452z2)) ;
    NAND3C NOT_FIFO_DEV_ix1455z50932 (.Y (nx1455z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx36356z2), .C (nx2452z2)) ;
    NAND3C NOT_FIFO_DEV_ix458z50932 (.Y (nx458z1), .A (NOT_FIFO_DEV_rtlc5n43_int
           ), .B (nx35359z2), .C (nx2452z2)) ;
    NAND3C NOT_FIFO_DEV_ix64997z50932 (.Y (nx64997z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx34362z2), .C (nx2452z2)) ;
    NAND3C NOT_FIFO_DEV_ix63001z50932 (.Y (nx63001z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx33365z2), .C (nx2452z2)) ;
    NAND3C NOT_FIFO_DEV_ix62004z50932 (.Y (nx62004z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx32368z2), .C (nx2452z2)) ;
    NAND3C NOT_FIFO_DEV_ix61007z50932 (.Y (nx61007z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx30372z2), .C (nx2452z2)) ;
    NAND3C NOT_FIFO_DEV_ix60010z50932 (.Y (nx60010z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx29375z2), .C (nx2452z2)) ;
    NAND3C NOT_FIFO_DEV_ix59013z50932 (.Y (nx59013z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx28378z2), .C (nx2452z2)) ;
    NAND3C NOT_FIFO_DEV_ix58016z50932 (.Y (nx58016z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx27381z2), .C (nx2452z2)) ;
    NAND3C NOT_FIFO_DEV_ix57019z50932 (.Y (nx57019z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx26384z2), .C (nx2452z2)) ;
    NAND3C NOT_FIFO_DEV_ix56022z50932 (.Y (nx56022z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx25387z2), .C (nx2452z2)) ;
    NAND3C NOT_FIFO_DEV_ix55025z50932 (.Y (nx55025z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx2452z2), .C (nx24390z2)) ;
    NAND3C NOT_FIFO_DEV_ix54028z50932 (.Y (nx54028z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx2452z2), .C (nx23393z2)) ;
    NAND3C NOT_FIFO_DEV_ix52032z50932 (.Y (nx52032z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx2452z2), .C (nx22396z2)) ;
    NAND3C NOT_FIFO_DEV_ix51035z50932 (.Y (nx51035z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx2452z2), .C (nx21399z2)) ;
    NAND3C NOT_FIFO_DEV_ix50038z50932 (.Y (nx50038z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx50038z2), .C (nx37353z4)) ;
    NAND3C NOT_FIFO_DEV_ix49041z50932 (.Y (nx49041z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx50038z2), .C (nx36356z2)) ;
    NAND3C NOT_FIFO_DEV_ix48044z50932 (.Y (nx48044z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx50038z2), .C (nx35359z2)) ;
    NAND3C NOT_FIFO_DEV_ix47047z50932 (.Y (nx47047z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx50038z2), .C (nx34362z2)) ;
    NAND3C NOT_FIFO_DEV_ix46050z50932 (.Y (nx46050z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx50038z2), .C (nx33365z2)) ;
    NAND3C NOT_FIFO_DEV_ix45053z50932 (.Y (nx45053z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx50038z2), .C (nx32368z2)) ;
    NAND3C NOT_FIFO_DEV_ix44056z50932 (.Y (nx44056z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx50038z2), .C (nx30372z2)) ;
    NAND3C NOT_FIFO_DEV_ix43059z50932 (.Y (nx43059z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx50038z2), .C (nx29375z2)) ;
    NAND3C NOT_FIFO_DEV_ix37436z50932 (.Y (nx37436z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx50038z2), .C (nx28378z2)) ;
    NAND3C NOT_FIFO_DEV_ix38433z50932 (.Y (nx38433z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx50038z2), .C (nx27381z2)) ;
    NAND3C NOT_FIFO_DEV_ix39430z50932 (.Y (nx39430z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx50038z2), .C (nx26384z2)) ;
    NAND3C NOT_FIFO_DEV_ix40427z50932 (.Y (nx40427z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx50038z2), .C (nx25387z2)) ;
    NAND3C NOT_FIFO_DEV_ix41424z50932 (.Y (nx41424z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx24390z2), .C (nx50038z2)) ;
    NAND3C NOT_FIFO_DEV_ix42421z50932 (.Y (nx42421z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx23393z2), .C (nx50038z2)) ;
    NAND3C NOT_FIFO_DEV_ix43418z50932 (.Y (nx43418z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx22396z2), .C (nx50038z2)) ;
    NAND3C NOT_FIFO_DEV_ix44415z50932 (.Y (nx44415z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx21399z2), .C (nx50038z2)) ;
    NAND3C NOT_FIFO_DEV_ix45412z50932 (.Y (nx45412z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx37353z4), .C (nx45412z2)) ;
    NAND3C NOT_FIFO_DEV_ix46409z50932 (.Y (nx46409z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx36356z2), .C (nx45412z2)) ;
    NAND3C NOT_FIFO_DEV_ix48405z50932 (.Y (nx48405z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx35359z2), .C (nx45412z2)) ;
    NAND3C NOT_FIFO_DEV_ix49402z50932 (.Y (nx49402z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx34362z2), .C (nx45412z2)) ;
    NAND3C NOT_FIFO_DEV_ix50399z50932 (.Y (nx50399z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx33365z2), .C (nx45412z2)) ;
    NAND3C NOT_FIFO_DEV_ix51396z50932 (.Y (nx51396z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx32368z2), .C (nx45412z2)) ;
    NAND3C NOT_FIFO_DEV_ix52393z50932 (.Y (nx52393z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx30372z2), .C (nx45412z2)) ;
    NAND3C NOT_FIFO_DEV_ix53390z50932 (.Y (nx53390z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx29375z2), .C (nx45412z2)) ;
    NAND3C NOT_FIFO_DEV_ix54387z50932 (.Y (nx54387z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx28378z2), .C (nx45412z2)) ;
    NAND3C NOT_FIFO_DEV_ix55384z50932 (.Y (nx55384z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx27381z2), .C (nx45412z2)) ;
    NAND3C NOT_FIFO_DEV_ix56381z50932 (.Y (nx56381z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx26384z2), .C (nx45412z2)) ;
    NAND3C NOT_FIFO_DEV_ix57378z50932 (.Y (nx57378z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx25387z2), .C (nx45412z2)) ;
    NAND3C NOT_FIFO_DEV_ix59374z50932 (.Y (nx59374z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx24390z2), .C (nx45412z2)) ;
    NAND3C NOT_FIFO_DEV_ix60371z50932 (.Y (nx60371z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx23393z2), .C (nx45412z2)) ;
    NAND3C NOT_FIFO_DEV_ix61368z50932 (.Y (nx61368z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx22396z2), .C (nx45412z2)) ;
    NAND3C NOT_FIFO_DEV_ix62365z50932 (.Y (nx62365z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx21399z2), .C (nx45412z2)) ;
    NAND3C NOT_FIFO_DEV_ix63362z50932 (.Y (nx63362z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx37353z4), .C (nx63362z2)) ;
    NAND3C NOT_FIFO_DEV_ix64359z50932 (.Y (nx64359z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx36356z2), .C (nx63362z2)) ;
    NAND3C NOT_FIFO_DEV_ix65356z50932 (.Y (nx65356z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx35359z2), .C (nx63362z2)) ;
    NAND3C NOT_FIFO_DEV_ix817z50932 (.Y (nx817z1), .A (NOT_FIFO_DEV_rtlc5n43_int
           ), .B (nx34362z2), .C (nx63362z2)) ;
    NAND3C NOT_FIFO_DEV_ix1814z50932 (.Y (nx1814z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx33365z2), .C (nx63362z2)) ;
    NAND3C NOT_FIFO_DEV_ix2811z50932 (.Y (nx2811z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx32368z2), .C (nx63362z2)) ;
    NAND3C NOT_FIFO_DEV_ix4807z50932 (.Y (nx4807z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx30372z2), .C (nx63362z2)) ;
    NAND3C NOT_FIFO_DEV_ix5804z50932 (.Y (nx5804z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx29375z2), .C (nx63362z2)) ;
    NAND3C NOT_FIFO_DEV_ix6801z50932 (.Y (nx6801z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx28378z2), .C (nx63362z2)) ;
    NAND3C NOT_FIFO_DEV_ix7798z50932 (.Y (nx7798z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx27381z2), .C (nx63362z2)) ;
    NAND3C NOT_FIFO_DEV_ix8795z50932 (.Y (nx8795z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx26384z2), .C (nx63362z2)) ;
    NAND3C NOT_FIFO_DEV_ix9792z50932 (.Y (nx9792z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx25387z2), .C (nx63362z2)) ;
    NAND3C NOT_FIFO_DEV_ix10789z50932 (.Y (nx10789z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx24390z2), .C (nx63362z2)) ;
    NAND3C NOT_FIFO_DEV_ix11786z50932 (.Y (nx11786z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx23393z2), .C (nx63362z2)) ;
    NAND3C NOT_FIFO_DEV_ix12783z50932 (.Y (nx12783z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx22396z2), .C (nx63362z2)) ;
    NAND3C NOT_FIFO_DEV_ix13780z50932 (.Y (nx13780z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx21399z2), .C (nx63362z2)) ;
    NAND3C NOT_FIFO_DEV_ix15776z50932 (.Y (nx15776z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx37353z4), .C (nx15776z2)) ;
    NAND3C NOT_FIFO_DEV_ix16773z50932 (.Y (nx16773z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx36356z2), .C (nx15776z2)) ;
    NAND3C NOT_FIFO_DEV_ix17770z50932 (.Y (nx17770z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx35359z2), .C (nx15776z2)) ;
    NAND3C NOT_FIFO_DEV_ix18767z50932 (.Y (nx18767z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx34362z2), .C (nx15776z2)) ;
    NAND3C NOT_FIFO_DEV_ix19764z50932 (.Y (nx19764z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx33365z2), .C (nx15776z2)) ;
    NAND3C NOT_FIFO_DEV_ix20761z50932 (.Y (nx20761z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx32368z2), .C (nx15776z2)) ;
    NAND3C NOT_FIFO_DEV_ix21758z50932 (.Y (nx21758z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx30372z2), .C (nx15776z2)) ;
    NAND3C NOT_FIFO_DEV_ix22755z50932 (.Y (nx22755z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx29375z2), .C (nx15776z2)) ;
    NAND3C NOT_FIFO_DEV_ix23752z50932 (.Y (nx23752z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx28378z2), .C (nx15776z2)) ;
    NAND3C NOT_FIFO_DEV_ix24749z50932 (.Y (nx24749z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx27381z2), .C (nx15776z2)) ;
    NAND3C NOT_FIFO_DEV_ix26745z50932 (.Y (nx26745z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx26384z2), .C (nx15776z2)) ;
    NAND3C NOT_FIFO_DEV_ix27742z50932 (.Y (nx27742z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx25387z2), .C (nx15776z2)) ;
    NAND3C NOT_FIFO_DEV_ix28739z50932 (.Y (nx28739z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx24390z2), .C (nx15776z2)) ;
    NAND3C NOT_FIFO_DEV_ix29736z50932 (.Y (nx29736z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx23393z2), .C (nx15776z2)) ;
    NAND3C NOT_FIFO_DEV_ix30733z50932 (.Y (nx30733z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx22396z2), .C (nx15776z2)) ;
    NAND3C NOT_FIFO_DEV_ix31730z50932 (.Y (nx31730z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx21399z2), .C (nx15776z2)) ;
    NAND3C NOT_FIFO_DEV_ix32727z50932 (.Y (nx32727z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx37353z4), .C (nx32727z2)) ;
    NAND3C NOT_FIFO_DEV_ix33724z50932 (.Y (nx33724z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx36356z2), .C (nx32727z2)) ;
    NAND3C NOT_FIFO_DEV_ix34721z50932 (.Y (nx34721z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx35359z2), .C (nx32727z2)) ;
    NAND3C NOT_FIFO_DEV_ix35718z50932 (.Y (nx35718z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx34362z2), .C (nx32727z2)) ;
    NAND3C NOT_FIFO_DEV_ix37714z50932 (.Y (nx37714z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx33365z2), .C (nx32727z2)) ;
    NAND3C NOT_FIFO_DEV_ix38711z50932 (.Y (nx38711z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx32368z2), .C (nx32727z2)) ;
    NAND3C NOT_FIFO_DEV_ix39708z50932 (.Y (nx39708z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx30372z2), .C (nx32727z2)) ;
    NAND3C NOT_FIFO_DEV_ix40705z50932 (.Y (nx40705z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx29375z2), .C (nx32727z2)) ;
    NAND3C NOT_FIFO_DEV_ix41702z50932 (.Y (nx41702z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx28378z2), .C (nx32727z2)) ;
    NAND3C NOT_FIFO_DEV_ix42699z50932 (.Y (nx42699z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx27381z2), .C (nx32727z2)) ;
    NAND3C NOT_FIFO_DEV_ix43696z50932 (.Y (nx43696z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx26384z2), .C (nx32727z2)) ;
    NAND3C NOT_FIFO_DEV_ix44693z50932 (.Y (nx44693z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx25387z2), .C (nx32727z2)) ;
    NAND3C NOT_FIFO_DEV_ix45690z50932 (.Y (nx45690z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx24390z2), .C (nx32727z2)) ;
    NAND3C NOT_FIFO_DEV_ix46687z50932 (.Y (nx46687z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx23393z2), .C (nx32727z2)) ;
    NAND3C NOT_FIFO_DEV_ix48683z50932 (.Y (nx48683z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx22396z2), .C (nx32727z2)) ;
    NAND3C NOT_FIFO_DEV_ix49680z50932 (.Y (nx49680z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx21399z2), .C (nx32727z2)) ;
    NAND3C NOT_FIFO_DEV_ix50677z50932 (.Y (nx50677z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx37353z4), .C (nx50677z2)) ;
    NAND3C NOT_FIFO_DEV_ix51674z50932 (.Y (nx51674z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx36356z2), .C (nx50677z2)) ;
    NAND3C NOT_FIFO_DEV_ix52671z50932 (.Y (nx52671z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx35359z2), .C (nx50677z2)) ;
    NAND3C NOT_FIFO_DEV_ix53668z50932 (.Y (nx53668z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx34362z2), .C (nx50677z2)) ;
    NAND3C NOT_FIFO_DEV_ix54665z50932 (.Y (nx54665z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx33365z2), .C (nx50677z2)) ;
    NAND3C NOT_FIFO_DEV_ix55662z50932 (.Y (nx55662z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx32368z2), .C (nx50677z2)) ;
    NAND3C NOT_FIFO_DEV_ix56659z50932 (.Y (nx56659z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx30372z2), .C (nx50677z2)) ;
    NAND3C NOT_FIFO_DEV_ix57656z50932 (.Y (nx57656z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx29375z2), .C (nx50677z2)) ;
    NAND3C NOT_FIFO_DEV_ix59652z50932 (.Y (nx59652z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx28378z2), .C (nx50677z2)) ;
    NAND3C NOT_FIFO_DEV_ix60649z50932 (.Y (nx60649z1), .A (nx50677z2), .B (
           nx27381z2), .C (NOT_FIFO_DEV_rtlc5n43_int)) ;
    NAND3C NOT_FIFO_DEV_ix61646z50932 (.Y (nx61646z1), .A (nx50677z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx26384z2)) ;
    NAND3C NOT_FIFO_DEV_ix62643z50932 (.Y (nx62643z1), .A (nx50677z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx25387z2)) ;
    NAND3C NOT_FIFO_DEV_ix63640z50932 (.Y (nx63640z1), .A (nx50677z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx24390z2)) ;
    NAND3C NOT_FIFO_DEV_ix64637z50932 (.Y (nx64637z1), .A (nx50677z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx23393z2)) ;
    NAND3C NOT_FIFO_DEV_ix98z50932 (.Y (nx98z1), .A (nx50677z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx22396z2)) ;
    NAND3C NOT_FIFO_DEV_ix1095z50932 (.Y (nx1095z1), .A (nx50677z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx21399z2)) ;
    NAND3C NOT_FIFO_DEV_ix2092z50932 (.Y (nx2092z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx2092z2), .C (nx37353z4)) ;
    NAND3C NOT_FIFO_DEV_ix3089z50932 (.Y (nx3089z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx2092z2), .C (nx36356z2)) ;
    NAND3C NOT_FIFO_DEV_ix5085z50932 (.Y (nx5085z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx2092z2), .C (nx35359z2)) ;
    NAND3C NOT_FIFO_DEV_ix6082z50932 (.Y (nx6082z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx2092z2), .C (nx34362z2)) ;
    NAND3C NOT_FIFO_DEV_ix7079z50932 (.Y (nx7079z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx2092z2), .C (nx33365z2)) ;
    NAND3C NOT_FIFO_DEV_ix8076z50932 (.Y (nx8076z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx2092z2), .C (nx32368z2)) ;
    NAND3C NOT_FIFO_DEV_ix9073z50932 (.Y (nx9073z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx2092z2), .C (nx30372z2)) ;
    NAND3C NOT_FIFO_DEV_ix10070z50932 (.Y (nx10070z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx2092z2), .C (nx29375z2)) ;
    NAND3C NOT_FIFO_DEV_ix11067z50932 (.Y (nx11067z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx2092z2), .C (nx28378z2)) ;
    NAND3C NOT_FIFO_DEV_ix12064z50932 (.Y (nx12064z1), .A (nx27381z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx2092z2)) ;
    NAND3C NOT_FIFO_DEV_ix13061z50932 (.Y (nx13061z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx26384z2), .C (nx2092z2)) ;
    NAND3C NOT_FIFO_DEV_ix14058z50932 (.Y (nx14058z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx25387z2), .C (nx2092z2)) ;
    NAND3C NOT_FIFO_DEV_ix5577z50932 (.Y (nx5577z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx24390z2), .C (nx2092z2)) ;
    NAND3C NOT_FIFO_DEV_ix6574z50932 (.Y (nx6574z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx23393z2), .C (nx2092z2)) ;
    NAND3C NOT_FIFO_DEV_ix7571z50932 (.Y (nx7571z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx22396z2), .C (nx2092z2)) ;
    NAND3C NOT_FIFO_DEV_ix8568z50932 (.Y (nx8568z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx21399z2), .C (nx2092z2)) ;
    NAND3C NOT_FIFO_DEV_ix9565z50932 (.Y (nx9565z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx37353z4), .C (nx9565z2)) ;
    NAND3C NOT_FIFO_DEV_ix10562z50932 (.Y (nx10562z4), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx36356z2), .C (nx9565z2)) ;
    NAND3C NOT_FIFO_DEV_ix11559z50932 (.Y (nx11559z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx35359z2), .C (nx9565z2)) ;
    NAND3C NOT_FIFO_DEV_ix12556z50932 (.Y (nx12556z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx34362z2), .C (nx9565z2)) ;
    NAND3C NOT_FIFO_DEV_ix13553z50932 (.Y (nx13553z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx33365z2), .C (nx9565z2)) ;
    NAND3C NOT_FIFO_DEV_ix14550z50932 (.Y (nx14550z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx32368z2), .C (nx9565z2)) ;
    NAND3C NOT_FIFO_DEV_ix16546z50932 (.Y (nx16546z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx30372z2), .C (nx9565z2)) ;
    NAND3C NOT_FIFO_DEV_ix17543z50932 (.Y (nx17543z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx29375z2), .C (nx9565z2)) ;
    NAND3C NOT_FIFO_DEV_ix18540z50932 (.Y (nx18540z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx28378z2), .C (nx9565z2)) ;
    NAND3C NOT_FIFO_DEV_ix19537z50932 (.Y (nx19537z1), .A (nx27381z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx9565z2)) ;
    NAND3C NOT_FIFO_DEV_ix20534z50932 (.Y (nx20534z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx26384z2), .C (nx9565z2)) ;
    NAND3C NOT_FIFO_DEV_ix21531z50932 (.Y (nx21531z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx25387z2), .C (nx9565z2)) ;
    NAND3C NOT_FIFO_DEV_ix22528z50932 (.Y (nx22528z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx24390z2), .C (nx9565z2)) ;
    NAND3C NOT_FIFO_DEV_ix23525z50932 (.Y (nx23525z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx23393z2), .C (nx9565z2)) ;
    NAND3C NOT_FIFO_DEV_ix24522z50932 (.Y (nx24522z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx22396z2), .C (nx9565z2)) ;
    NAND3C NOT_FIFO_DEV_ix25519z50932 (.Y (nx25519z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx21399z2), .C (nx9565z2)) ;
    NAND3C NOT_FIFO_DEV_ix27515z50932 (.Y (nx27515z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx37353z4), .C (nx27515z2)) ;
    NAND3C NOT_FIFO_DEV_ix28512z50932 (.Y (nx28512z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx36356z2), .C (nx27515z2)) ;
    NAND3C NOT_FIFO_DEV_ix29509z50932 (.Y (nx29509z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx35359z2), .C (nx27515z2)) ;
    NAND3C NOT_FIFO_DEV_ix30506z50932 (.Y (nx30506z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx34362z2), .C (nx27515z2)) ;
    NAND3C NOT_FIFO_DEV_ix31503z50932 (.Y (nx31503z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx33365z2), .C (nx27515z2)) ;
    NAND3C NOT_FIFO_DEV_ix32500z50932 (.Y (nx32500z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx32368z2), .C (nx27515z2)) ;
    NAND3C NOT_FIFO_DEV_ix33497z50932 (.Y (nx33497z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx30372z2), .C (nx27515z2)) ;
    NAND3C NOT_FIFO_DEV_ix34494z50932 (.Y (nx34494z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx29375z2), .C (nx27515z2)) ;
    NAND3C NOT_FIFO_DEV_ix35491z50932 (.Y (nx35491z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx28378z2), .C (nx27515z2)) ;
    NAND3C NOT_FIFO_DEV_ix36488z50932 (.Y (nx36488z1), .A (nx27381z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx27515z2)) ;
    NAND3C NOT_FIFO_DEV_ix38484z50932 (.Y (nx38484z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx26384z2), .C (nx27515z2)) ;
    NAND3C NOT_FIFO_DEV_ix39481z50932 (.Y (nx39481z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx25387z2), .C (nx27515z2)) ;
    NAND3C NOT_FIFO_DEV_ix40478z50932 (.Y (nx40478z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx24390z2), .C (nx27515z2)) ;
    NAND3C NOT_FIFO_DEV_ix41475z50932 (.Y (nx41475z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx23393z2), .C (nx27515z2)) ;
    NAND3C NOT_FIFO_DEV_ix42472z50932 (.Y (nx42472z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx22396z2), .C (nx27515z2)) ;
    NAND3C NOT_FIFO_DEV_ix43469z50932 (.Y (nx43469z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx21399z2), .C (nx27515z2)) ;
    NAND3C NOT_FIFO_DEV_ix44466z50932 (.Y (nx44466z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx37353z4), .C (nx44466z2)) ;
    NAND3C NOT_FIFO_DEV_ix45463z50932 (.Y (nx45463z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx36356z2), .C (nx44466z2)) ;
    NAND3C NOT_FIFO_DEV_ix46460z50932 (.Y (nx46460z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx35359z2), .C (nx44466z2)) ;
    NAND3C NOT_FIFO_DEV_ix47457z50932 (.Y (nx47457z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx34362z2), .C (nx44466z2)) ;
    NAND3C NOT_FIFO_DEV_ix49453z50932 (.Y (nx49453z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx33365z2), .C (nx44466z2)) ;
    NAND3C NOT_FIFO_DEV_ix50450z50932 (.Y (nx50450z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx32368z2), .C (nx44466z2)) ;
    NAND3C NOT_FIFO_DEV_ix51447z50932 (.Y (nx51447z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx30372z2), .C (nx44466z2)) ;
    NAND3C NOT_FIFO_DEV_ix52444z50932 (.Y (nx52444z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx29375z2), .C (nx44466z2)) ;
    NAND3C NOT_FIFO_DEV_ix53441z50932 (.Y (nx53441z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx28378z2), .C (nx44466z2)) ;
    NAND3C NOT_FIFO_DEV_ix54438z50932 (.Y (nx54438z1), .A (nx27381z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx44466z2)) ;
    NAND3C NOT_FIFO_DEV_ix55435z50932 (.Y (nx55435z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx26384z2), .C (nx44466z2)) ;
    NAND3C NOT_FIFO_DEV_ix56432z50932 (.Y (nx56432z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx25387z2), .C (nx44466z2)) ;
    NAND3C NOT_FIFO_DEV_ix57429z50932 (.Y (nx57429z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx24390z2), .C (nx44466z2)) ;
    NAND3C NOT_FIFO_DEV_ix58426z50932 (.Y (nx58426z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx23393z2), .C (nx44466z2)) ;
    NAND3C NOT_FIFO_DEV_ix60422z50932 (.Y (nx60422z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx22396z2), .C (nx44466z2)) ;
    NAND3C NOT_FIFO_DEV_ix61419z50932 (.Y (nx61419z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx21399z2), .C (nx44466z2)) ;
    NAND3C NOT_FIFO_DEV_ix62416z50932 (.Y (nx62416z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx37353z4), .C (nx62416z2)) ;
    NAND3C NOT_FIFO_DEV_ix63413z50932 (.Y (nx63413z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx36356z2), .C (nx62416z2)) ;
    NAND3C NOT_FIFO_DEV_ix64410z50932 (.Y (nx64410z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx35359z2), .C (nx62416z2)) ;
    NAND3C NOT_FIFO_DEV_ix65407z50932 (.Y (nx65407z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx34362z2), .C (nx62416z2)) ;
    NAND3C NOT_FIFO_DEV_ix868z50932 (.Y (nx868z1), .A (NOT_FIFO_DEV_rtlc5n43_int
           ), .B (nx33365z2), .C (nx62416z2)) ;
    NAND3C NOT_FIFO_DEV_ix1865z50932 (.Y (nx1865z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx32368z2), .C (nx62416z2)) ;
    NAND3C NOT_FIFO_DEV_ix2862z50932 (.Y (nx2862z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx30372z2), .C (nx62416z2)) ;
    NAND3C NOT_FIFO_DEV_ix3859z50932 (.Y (nx3859z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx29375z2), .C (nx62416z2)) ;
    NAND3C NOT_FIFO_DEV_ix5855z50932 (.Y (nx5855z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx28378z2), .C (nx62416z2)) ;
    NAND3C NOT_FIFO_DEV_ix6852z50932 (.Y (nx6852z1), .A (nx27381z2), .B (
           NOT_FIFO_DEV_rtlc5n43_int), .C (nx62416z2)) ;
    NAND3C NOT_FIFO_DEV_ix7849z50932 (.Y (nx7849z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx26384z2), .C (nx62416z2)) ;
    NAND3C NOT_FIFO_DEV_ix8846z50932 (.Y (nx8846z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx25387z2), .C (nx62416z2)) ;
    NAND3C NOT_FIFO_DEV_ix9843z50932 (.Y (nx9843z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx24390z2), .C (nx62416z2)) ;
    NAND3C NOT_FIFO_DEV_ix10840z50932 (.Y (nx10840z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx23393z2), .C (nx62416z2)) ;
    NAND3C NOT_FIFO_DEV_ix11837z50932 (.Y (nx11837z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx22396z2), .C (nx62416z2)) ;
    NAND3C NOT_FIFO_DEV_ix12834z50932 (.Y (nx12834z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx21399z2), .C (nx62416z2)) ;
    NAND3C NOT_FIFO_DEV_ix13831z50932 (.Y (nx13831z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx37353z4), .C (nx13831z2)) ;
    NAND3C NOT_FIFO_DEV_ix14828z50932 (.Y (nx14828z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx36356z2), .C (nx13831z2)) ;
    NAND3C NOT_FIFO_DEV_ix16824z50932 (.Y (nx16824z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx35359z2), .C (nx13831z2)) ;
    NAND3C NOT_FIFO_DEV_ix17821z50932 (.Y (nx17821z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx34362z2), .C (nx13831z2)) ;
    NAND3C NOT_FIFO_DEV_ix18818z50932 (.Y (nx18818z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx33365z2), .C (nx13831z2)) ;
    NAND3C NOT_FIFO_DEV_ix19815z50932 (.Y (nx19815z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx32368z2), .C (nx13831z2)) ;
    NAND3C NOT_FIFO_DEV_ix20812z50932 (.Y (nx20812z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx13831z2), .C (nx30372z2)) ;
    NAND3C NOT_FIFO_DEV_ix21809z50932 (.Y (nx21809z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx13831z2), .C (nx29375z2)) ;
    NAND3C NOT_FIFO_DEV_ix22806z50932 (.Y (nx22806z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx13831z2), .C (nx28378z2)) ;
    NAND3C NOT_FIFO_DEV_ix23803z50932 (.Y (nx23803z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx13831z2), .C (nx27381z2)) ;
    NAND3C NOT_FIFO_DEV_ix24800z50932 (.Y (nx24800z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx13831z2), .C (nx26384z2)) ;
    NAND3C NOT_FIFO_DEV_ix25797z50932 (.Y (nx25797z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx13831z2), .C (nx25387z2)) ;
    NAND3C NOT_FIFO_DEV_ix27793z50932 (.Y (nx27793z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx13831z2), .C (nx24390z2)) ;
    NAND3C NOT_FIFO_DEV_ix28790z50932 (.Y (nx28790z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx13831z2), .C (nx23393z2)) ;
    NAND3C NOT_FIFO_DEV_ix29787z50932 (.Y (nx29787z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx13831z2), .C (nx22396z2)) ;
    NAND3C NOT_FIFO_DEV_ix30784z50932 (.Y (nx30784z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx13831z2), .C (nx21399z2)) ;
    NAND3C NOT_FIFO_DEV_ix31781z50932 (.Y (nx31781z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx31781z2), .C (nx37353z4)) ;
    NAND3C NOT_FIFO_DEV_ix32778z50932 (.Y (nx32778z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx31781z2), .C (nx36356z2)) ;
    NAND3C NOT_FIFO_DEV_ix33775z50932 (.Y (nx33775z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx31781z2), .C (nx35359z2)) ;
    NAND3C NOT_FIFO_DEV_ix34772z50932 (.Y (nx34772z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx31781z2), .C (nx34362z2)) ;
    NAND3C NOT_FIFO_DEV_ix35769z50932 (.Y (nx35769z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx31781z2), .C (nx33365z2)) ;
    NAND3C NOT_FIFO_DEV_ix36766z50932 (.Y (nx36766z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx32368z2), .C (nx31781z2)) ;
    NAND3C NOT_FIFO_DEV_ix48358z50932 (.Y (nx48358z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx30372z2), .C (nx31781z2)) ;
    NAND3C NOT_FIFO_DEV_ix47361z50932 (.Y (nx47361z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx29375z2), .C (nx31781z2)) ;
    NAND3C NOT_FIFO_DEV_ix46364z50932 (.Y (nx46364z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx28378z2), .C (nx31781z2)) ;
    NAND3C NOT_FIFO_DEV_ix45367z50932 (.Y (nx45367z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx27381z2), .C (nx31781z2)) ;
    NAND3C NOT_FIFO_DEV_ix44370z50932 (.Y (nx44370z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx26384z2), .C (nx31781z2)) ;
    NAND3C NOT_FIFO_DEV_ix43373z50932 (.Y (nx43373z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx25387z2), .C (nx31781z2)) ;
    NAND3C NOT_FIFO_DEV_ix42376z50932 (.Y (nx42376z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx24390z2), .C (nx31781z2)) ;
    NAND3C NOT_FIFO_DEV_ix41379z50932 (.Y (nx41379z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx23393z2), .C (nx31781z2)) ;
    NAND3C NOT_FIFO_DEV_ix40382z50932 (.Y (nx40382z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx22396z2), .C (nx31781z2)) ;
    NAND3C NOT_FIFO_DEV_ix39385z50932 (.Y (nx39385z1), .A (
           NOT_FIFO_DEV_rtlc5n43_int), .B (nx21399z2), .C (nx31781z2)) ;
    NAND2 ix12521z24339 (.Y (nx12521z2), .A (CONDITION_1_), .B (READ_int)) ;
    XO1A FIFO_DEV_rtlc14_X_0_n123_rename1014 (.Y (FIFO_DEV_rtlc14_X_0_n123), .A (
         WRITE), .B (READ_int), .C (nx59980z1)) ;
    AO1E NOT_ENCR_DEV_modgen_counter_key_cnt_ix45632z40560 (.Y (nx45632z2), .A (
         ENCR_DEV_rtlc12_X_0_n169), .B (ENCR_DEV_prev_1___repl0), .C (nx45632z3)
         ) ;
    XO1A ix22484z43526 (.Y (nx22484z1), .A (NOT_ENCR_DEV_t_1_4_16n1s20), .B (
         nx22484z2), .C (NOT_ENCR_DEV_rtlcn261_int)) ;
    XO1A ix25475z43526 (.Y (nx25475z1), .A (NOT_ENCR_DEV_t_1_7_16n1s32), .B (
         nx25475z2), .C (NOT_ENCR_DEV_rtlcn261_int)) ;
    NAND3 ix5542z24339 (.Y (nx5542z3), .A (nx12521z4), .B (nx12521z8), .C (
          nx5542z4)) ;
    NAND3 ix6539z24339 (.Y (nx6539z3), .A (nx12521z4), .B (nx12521z8), .C (
          nx6539z4)) ;
    NAND3 ix7536z24339 (.Y (nx7536z3), .A (nx12521z4), .B (nx12521z8), .C (
          nx7536z4)) ;
    NAND3 ix8533z24339 (.Y (nx8533z3), .A (nx12521z4), .B (nx12521z8), .C (
          nx8533z4)) ;
    NAND3 ix9530z24339 (.Y (nx9530z3), .A (nx12521z4), .B (nx12521z8), .C (
          nx9530z4)) ;
    NAND3 ix10527z24339 (.Y (nx10527z3), .A (nx12521z4), .B (nx12521z8), .C (
          nx10527z4)) ;
    NAND3 ix11524z24339 (.Y (nx11524z3), .A (nx12521z4), .B (nx12521z8), .C (
          nx11524z4)) ;
    NAND3 ix12521z24343 (.Y (nx12521z7), .A (nx12521z4), .B (nx12521z8), .C (
          nx12521z11)) ;
    NAND3A ix35840z50931 (.Y (nx35840z2), .A (b_0__int), .B (
           NOT_ENCR_DEV_rtlcn261_int), .C (ENCR_DEV_key_reg[2])) ;
    NAND3A ix42819z50931 (.Y (nx42819z2), .A (b_0__int), .B (
           NOT_ENCR_DEV_rtlcn261_int), .C (ENCR_DEV_key_reg[9])) ;
    NAND3A ix25475z50932 (.Y (nx25475z3), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
           b_0__int), .C (ENCR_DEV_t_1_0_)) ;
    NAND3A ix22484z50932 (.Y (nx22484z3), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
           b_0__int), .C (ENCR_DEV_reg_str_2[2])) ;
    NAND2 ix17499z24338 (.Y (nx17499z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[7])) ;
    AO1D ix17499z40559 (.Y (nx17499z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[0]), .C (b_0__int)) ;
    NAND2 ix47382z24338 (.Y (nx47382z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[9])) ;
    AO1D ix47382z40559 (.Y (nx47382z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[2]), .C (b_0__int)) ;
    NAND2 ix50373z24338 (.Y (nx50373z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[12])) ;
    AO1D ix50373z40559 (.Y (nx50373z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[5]), .C (b_0__int)) ;
    NAND2 ix51370z24338 (.Y (nx51370z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[13])) ;
    AO1D ix51370z40559 (.Y (nx51370z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[6]), .C (b_0__int)) ;
    NAND2 ix54361z24338 (.Y (nx54361z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[16])) ;
    AO1D ix54361z40559 (.Y (nx54361z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[9]), .C (b_0__int)) ;
    NAND2 ix55358z24338 (.Y (nx55358z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[17])) ;
    AO1D ix55358z40559 (.Y (nx55358z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[10]), .C (b_0__int)) ;
    NAND2 ix60345z24338 (.Y (nx60345z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[21])) ;
    AO1D ix60345z40559 (.Y (nx60345z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[14]), .C (b_0__int)) ;
    NAND2 ix791z24338 (.Y (nx791z1), .A (b_0__int), .B (ENCR_DEV_reg_str_2[27])
          ) ;
    AO1D ix791z40559 (.Y (nx791z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[20]), .C (b_0__int)) ;
    NAND2 ix1788z24338 (.Y (nx1788z1), .A (b_0__int), .B (ENCR_DEV_reg_str_2[28]
          )) ;
    AO1D ix1788z40559 (.Y (nx1788z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[21]), .C (b_0__int)) ;
    NAND2 ix3784z24338 (.Y (nx3784z1), .A (b_0__int), .B (ENCR_DEV_reg_str_2[29]
          )) ;
    AO1D ix3784z40559 (.Y (nx3784z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[22]), .C (b_0__int)) ;
    NAND2 ix7772z24338 (.Y (nx7772z1), .A (b_0__int), .B (ENCR_DEV_reg_str_2[33]
          )) ;
    AO1D ix7772z40559 (.Y (nx7772z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[26]), .C (b_0__int)) ;
    NAND2 ix9766z24338 (.Y (nx9766z1), .A (b_0__int), .B (ENCR_DEV_reg_str_2[35]
          )) ;
    AO1D ix9766z40559 (.Y (nx9766z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[28]), .C (b_0__int)) ;
    NAND2 ix11760z24338 (.Y (nx11760z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[37])) ;
    AO1D ix11760z40559 (.Y (nx11760z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[30]), .C (b_0__int)) ;
    NAND2 ix12757z24338 (.Y (nx12757z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[38])) ;
    AO1D ix12757z40559 (.Y (nx12757z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[31]), .C (b_0__int)) ;
    NAND2 ix15750z24338 (.Y (nx15750z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[40])) ;
    AO1D ix15750z40559 (.Y (nx15750z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[33]), .C (b_0__int)) ;
    NAND2 ix16747z24338 (.Y (nx16747z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[41])) ;
    AO1D ix16747z40559 (.Y (nx16747z2), .A (ENCR_DEV_reg_str_2[34]), .B (
         NOT_ENCR_DEV_rtlcn261_int), .C (b_0__int)) ;
    NAND2 ix18741z24338 (.Y (nx18741z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[43])) ;
    AO1D ix18741z40559 (.Y (nx18741z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[36]), .C (b_0__int)) ;
    NAND2 ix20735z24338 (.Y (nx20735z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[45])) ;
    AO1D ix20735z40559 (.Y (nx20735z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[38]), .C (b_0__int)) ;
    NAND2 ix22729z24338 (.Y (nx22729z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[47])) ;
    AO1D ix22729z40559 (.Y (nx22729z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[40]), .C (b_0__int)) ;
    NAND2 ix23726z24338 (.Y (nx23726z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[48])) ;
    AO1D ix23726z40559 (.Y (nx23726z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[41]), .C (b_0__int)) ;
    NAND2 ix26719z24338 (.Y (nx26719z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[50])) ;
    AO1D ix26719z40559 (.Y (nx26719z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[43]), .C (b_0__int)) ;
    NAND2 ix27716z24338 (.Y (nx27716z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[51])) ;
    AO1D ix27716z40559 (.Y (nx27716z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[44]), .C (b_0__int)) ;
    NAND2 ix29710z24338 (.Y (nx29710z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[53])) ;
    AO1D ix29710z40559 (.Y (nx29710z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[46]), .C (b_0__int)) ;
    NAND2 ix31704z24338 (.Y (nx31704z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[55])) ;
    AO1D ix31704z40559 (.Y (nx31704z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[48]), .C (b_0__int)) ;
    NAND2 ix36691z24338 (.Y (nx36691z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[59])) ;
    AO1D ix36691z40559 (.Y (nx36691z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[52]), .C (b_0__int)) ;
    NAND2 ix37688z24340 (.Y (nx37688z2), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[60])) ;
    AO1D ix37688z40561 (.Y (nx37688z3), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[53]), .C (b_0__int)) ;
    NAND2 ix38685z24338 (.Y (nx38685z1), .A (ENCR_DEV_reg_str_2[61]), .B (
          b_0__int)) ;
    AO1D ix38685z40559 (.Y (nx38685z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[54]), .C (b_0__int)) ;
    NAND2 ix41676z24338 (.Y (nx41676z1), .A (ENCR_DEV_reg_str_2[64]), .B (
          b_0__int)) ;
    AO1D ix41676z40559 (.Y (nx41676z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[57]), .C (b_0__int)) ;
    NAND2 ix42673z24338 (.Y (nx42673z1), .A (ENCR_DEV_reg_str_2[65]), .B (
          b_0__int)) ;
    AO1D ix42673z40559 (.Y (nx42673z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[58]), .C (b_0__int)) ;
    NAND2 ix48657z24338 (.Y (nx48657z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_2[70])) ;
    AO1D ix48657z40559 (.Y (nx48657z2), .A (ENCR_DEV_reg_str_2[63]), .B (
         NOT_ENCR_DEV_rtlcn261_int), .C (b_0__int)) ;
    NAND2 ix50651z24338 (.Y (nx50651z1), .A (ENCR_DEV_reg_str_2[72]), .B (
          b_0__int)) ;
    AO1D ix50651z40559 (.Y (nx50651z2), .A (ENCR_DEV_reg_str_2[65]), .B (
         NOT_ENCR_DEV_rtlcn261_int), .C (b_0__int)) ;
    NAND2 ix51648z24338 (.Y (nx51648z1), .A (ENCR_DEV_reg_str_2[73]), .B (
          b_0__int)) ;
    AO1D ix51648z40559 (.Y (nx51648z2), .A (ENCR_DEV_reg_str_2[66]), .B (
         NOT_ENCR_DEV_rtlcn261_int), .C (b_0__int)) ;
    NAND2 ix55636z24338 (.Y (nx55636z1), .A (ENCR_DEV_reg_str_2[77]), .B (
          b_0__int)) ;
    AO1D ix55636z40559 (.Y (nx55636z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[70]), .C (b_0__int)) ;
    NAND2 ix56633z24338 (.Y (nx56633z1), .A (ENCR_DEV_reg_str_2[78]), .B (
          b_0__int)) ;
    AO1D ix56633z40559 (.Y (nx56633z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_2[71]), .C (b_0__int)) ;
    NAND2 ix35127z24338 (.Y (nx35127z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_3[107])) ;
    AO1D ix35127z40559 (.Y (nx35127z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_3[100]), .C (b_0__int)) ;
    NAND2 ix36124z24338 (.Y (nx36124z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_3[108])) ;
    AO1D ix36124z40559 (.Y (nx36124z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_3[101]), .C (b_0__int)) ;
    NAND2 ix38120z24338 (.Y (nx38120z1), .A (b_0__int), .B (
          ENCR_DEV_reg_str_3[109])) ;
    AO1D ix38120z40559 (.Y (nx38120z2), .A (NOT_ENCR_DEV_rtlcn261_int), .B (
         ENCR_DEV_reg_str_3[102]), .C (b_0__int)) ;
    NAND3B ix11504z50949 (.Y (nx11504z18), .A (STB_KEY_int), .B (nx11504z19), .C (
           ENCR_DEV_prev[2])) ;
    NAND3B ix65298z50931 (.Y (nx65298z1), .A (nx37353z3), .B (nx49948z1), .C (
           FIFO_DEV_rtlc_wadd_n4[6])) ;
    NAND3 ix32158z24340 (.Y (nx32158z3), .A (FIFO_DEV_rtlc_wadd_n4[4]), .B (
          FIFO_DEV_rtlc_wadd_n4[3]), .C (FIFO_DEV_rtlc_wadd_n4[2])) ;
    AND3B ix14495z2957 (.Y (nx14495z1), .A (STB_KEY_int), .B (nx14495z2), .C (
          ENCR_DEV_prev_1___repl0)) ;
    AND2 ix12521z48518 (.Y (nx12521z5), .A (CONDITION_1_), .B (READ_int)) ;
    MX2C ix12521z26299 (.Y (FIFO_DEV_not_dout_2n1s3), .A (nx12521z9), .S (
         FIFO_DEV_rtlc_radd_N1[7]), .B (nx12521z10)) ;
    NAND3C ix10562z50932 (.Y (nx10562z1), .A (nx10562z2), .B (nx6004z1), .C (
           nx31484z2)) ;
    NAND3C ix6418z50932 (.Y (nx6418z1), .A (nx6418z2), .B (nx14918z4), .C (
           nx19748z3)) ;
    NAND3C ix11504z50934 (.Y (NOT_a_7_), .A (nx11504z3), .B (nx49501z8), .C (
           nx8409z3)) ;
    NAND3C ix20284z50934 (.Y (NOT_a_1__dup_3637), .A (nx20284z3), .B (nx35506z5)
           , .C (nx55510z3)) ;
    NAND3C ix22498z50934 (.Y (NOT_a_1_), .A (nx22498z3), .B (nx52784z5), .C (
           nx52808z3)) ;
    NAND3C ix65280z50933 (.Y (NOT_a_1__dup_3625), .A (nx65280z2), .B (nx55534z4)
           , .C (nx35482z3)) ;
    NAND3A ix16808z50930 (.Y (nx16808z1), .A (nx49948z1), .B (
           FIFO_DEV_rtlc_wadd_n4[5]), .C (FIFO_DEV_rtlc_wadd_n4[4])) ;
    XOR2 ix10274z10876 (.Y (FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_1_), .A (
         FIFO_DEV_rtlc_radd_N1_0___repl0), .B (FIFO_DEV_rtlc_radd_N1_1___repl0)
         ) ;
    XOR2 ix48026z10877 (.Y (nx48026z2), .A (ENCR_DEV_reg_str_1[92]), .B (
         ENCR_DEV_reg_str_3[110])) ;
    XOR2 ix47029z10877 (.Y (nx47029z2), .A (ENCR_DEV_reg_str_3[64]), .B (
         ENCR_DEV_reg_str_2[67])) ;
    XOR2 ix46032z10877 (.Y (nx46032z2), .A (ENCR_DEV_reg_str_3[63]), .B (
         ENCR_DEV_reg_str_2[66])) ;
    XOR2 ix45035z10877 (.Y (nx45035z2), .A (ENCR_DEV_reg_str_3[62]), .B (
         ENCR_DEV_reg_str_2[65])) ;
    XOR2 ix44038z10877 (.Y (nx44038z2), .A (ENCR_DEV_reg_str_3[61]), .B (
         ENCR_DEV_reg_str_2[64])) ;
    XOR2 ix43041z10877 (.Y (nx43041z2), .A (ENCR_DEV_reg_str_2[63]), .B (
         ENCR_DEV_reg_str_3[60])) ;
    XOR2 ix42044z10877 (.Y (nx42044z2), .A (ENCR_DEV_reg_str_2[62]), .B (
         ENCR_DEV_reg_str_3[104])) ;
    XOR2 ix41047z10877 (.Y (nx41047z2), .A (ENCR_DEV_reg_str_2[61]), .B (
         ENCR_DEV_reg_str_3[58])) ;
    DFN1C0 ENCR_DEV_reg_sign_reg_4_ (.Q (SIGN_REG_dup_0[6]), .D (
           ENCR_DEV_prev_6__int), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_sign_reg_3_ (.Q (SIGN_REG_dup_0[5]), .D (
           ENCR_DEV_prev_5___repl0), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_sign_reg_2_ (.Q (SIGN_REG_dup_0[4]), .D (
           ENCR_DEV_prev[4]), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_sign_reg_1_ (.Q (SIGN_REG_dup_0[3]), .D (
           ENCR_DEV_prev[3]), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_sign_reg_0_ (.Q (SIGN_REG_dup_0[2]), .D (
           ENCR_DEV_prev[2]), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ix12521z38802 (.Q (nx12521z1), .D (ENCR_DEV_PWR), .E (nx12521z2), .CLK (
             CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_prev_6_ (.Q (ENCR_DEV_prev[6]), .D (nx13498z1), .CLK (
           CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_prev_5_ (.Q (ENCR_DEV_prev[5]), .D (nx36622z1), .CLK (
           CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_prev_4_ (.Q (ENCR_DEV_prev[4]), .D (nx11504z1), .CLK (
           CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_prev_3_ (.Q (ENCR_DEV_prev[3]), .D (nx10507z1), .CLK (
           CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_prev_2_ (.Q (ENCR_DEV_prev[2]), .D (nx9510z1), .CLK (
           CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_stream_7_ (.Q (STREAM[7]), .D (
             ENCR_DEV_stream_15n2ss1[7]), .E (nx46110z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_stream_6_ (.Q (STREAM[6]), .D (
             ENCR_DEV_stream_15n2ss1[6]), .E (nx46110z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_stream_5_ (.Q (STREAM[5]), .D (
             ENCR_DEV_stream_15n2ss1[5]), .E (nx46110z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_stream_4_ (.Q (STREAM[4]), .D (
             ENCR_DEV_stream_15n2ss1[4]), .E (nx46110z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_stream_3_ (.Q (STREAM[3]), .D (
             ENCR_DEV_stream_15n2ss1[3]), .E (nx46110z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_stream_2_ (.Q (STREAM[2]), .D (
             ENCR_DEV_stream_15n2ss1[2]), .E (nx46110z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_stream_1_ (.Q (STREAM[1]), .D (
             ENCR_DEV_stream_15n2ss1[1]), .E (nx46110z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_stream_0_ (.Q (STREAM[0]), .D (
             ENCR_DEV_stream_15n2ss1[0]), .E (nx46110z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1C0 reg_q_7__dup_42 (.Q (FIFO_DEV_rtlc_wadd_n4[7]), .D (inc_d_7__dup_2804
           ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 reg_q_6__dup_43 (.Q (FIFO_DEV_rtlc_wadd_n4[6]), .D (inc_d_6__dup_2803
           ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 reg_q_5__dup_44 (.Q (FIFO_DEV_rtlc_wadd_n4[5]), .D (inc_d_5__dup_2802
           ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 reg_q_4__dup_45 (.Q (FIFO_DEV_rtlc_wadd_n4[4]), .D (inc_d_4__dup_2801
           ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 reg_q_3__dup_46 (.Q (FIFO_DEV_rtlc_wadd_n4[3]), .D (inc_d_3__dup_2800
           ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 reg_q_2__dup_47 (.Q (FIFO_DEV_rtlc_wadd_n4[2]), .D (inc_d_2__dup_2799
           ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 reg_q_1__dup_48 (.Q (FIFO_DEV_rtlc_wadd_n4[1]), .D (inc_d_1__dup_2798
           ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 reg_q_0__dup_49 (.Q (FIFO_DEV_rtlc_wadd_n4[0]), .D (inc_d_0__dup_2797
           ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 FIFO_DEV_modgen_counter_rtlc_radd_N1_reg_q_7__dup (.Q (
             FIFO_DEV_rtlc_radd_N1[7]), .D (
             FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_7_), .E (nx12521z2), .CLK (
             CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 FIFO_DEV_modgen_counter_rtlc_radd_N1_reg_q_6__dup (.Q (
             FIFO_DEV_rtlc_radd_N1[6]), .D (
             FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_6_), .E (nx12521z2), .CLK (
             CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 FIFO_DEV_modgen_counter_rtlc_radd_N1_reg_q_5__dup (.Q (
             FIFO_DEV_rtlc_radd_N1[5]), .D (
             FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_5_), .E (nx12521z2), .CLK (
             CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 FIFO_DEV_modgen_counter_rtlc_radd_N1_reg_q_4__dup (.Q (
             FIFO_DEV_rtlc_radd_N1[4]), .D (
             FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_4_), .E (nx12521z2), .CLK (
             CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 FIFO_DEV_modgen_counter_rtlc_radd_N1_reg_q_3__dup (.Q (
             FIFO_DEV_rtlc_radd_N1[3]), .D (
             FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_3_), .E (nx12521z2), .CLK (
             CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 FIFO_DEV_modgen_counter_rtlc_radd_N1_reg_q_2__dup (.Q (
             FIFO_DEV_rtlc_radd_N1[2]), .D (
             FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_2_), .E (nx12521z2), .CLK (
             CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 FIFO_DEV_modgen_counter_rtlc_radd_N1_reg_q_1__dup (.Q (
             FIFO_DEV_rtlc_radd_N1[1]), .D (
             FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_1_), .E (nx12521z2), .CLK (
             CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 FIFO_DEV_modgen_counter_rtlc_radd_N1_reg_q_0__dup (.Q (
             FIFO_DEV_rtlc_radd_N1[0]), .D (
             FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_0_), .E (nx12521z2), .CLK (
             CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_wt_sgn (.Q (WRITE), .D (nx1908z1), .E (
             ENCR_DEV_rtlc15_PS14_n166), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_prev_1_ (.Q (ENCR_DEV_prev[1]), .D (nx3438z1), .CLK (
           CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_modgen_counter_key_cnt_reg_q_6_ (.Q (ENCR_DEV_key_cnt[6])
             , .D (nx39650z1), .E (nx45632z2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_prev_8_ (.Q (ENCR_DEV_prev[8]), .D (nx15492z1), .CLK (
           CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_5__dup_52 (.Q (FIFO_DEV_count[5]), .D (incdec_mux_5_dup_103)
             , .E (FIFO_DEV_rtlc14_X_0_n123), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_4__dup_53 (.Q (FIFO_DEV_count[4]), .D (incdec_mux_4_dup_102)
             , .E (FIFO_DEV_rtlc14_X_0_n123), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_3__dup_54 (.Q (FIFO_DEV_count[3]), .D (incdec_mux_3_dup_101)
             , .E (FIFO_DEV_rtlc14_X_0_n123), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_2__dup_55 (.Q (FIFO_DEV_count[2]), .D (incdec_mux_2_dup_100)
             , .E (FIFO_DEV_rtlc14_X_0_n123), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_1__dup_56 (.Q (FIFO_DEV_count[1]), .D (incdec_mux_1_dup_99), 
             .E (FIFO_DEV_rtlc14_X_0_n123), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_0__dup_57 (.Q (FIFO_DEV_count[0]), .D (a_0__dup_2819), .E (
             FIFO_DEV_rtlc14_X_0_n123), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_modgen_counter_key_cnt_reg_q_5_ (.Q (ENCR_DEV_key_cnt[5])
             , .D (nx40647z1), .E (nx45632z2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_modgen_counter_key_cnt_reg_q_4_ (.Q (ENCR_DEV_key_cnt[4])
             , .D (nx41644z1), .E (nx45632z2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_modgen_counter_key_cnt_reg_q_3_ (.Q (ENCR_DEV_key_cnt[3])
             , .D (nx42641z1), .E (nx45632z2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_modgen_counter_key_cnt_reg_q_2_ (.Q (ENCR_DEV_key_cnt[2])
             , .D (nx43638z1), .E (nx45632z2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_0__dup_32 (.Q (ENCR_DEV_encry_cnt[0]), .D (
             sclear_and_0_dup_114), .E (nx25368z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1C0 reg_q_11_ (.Q (ENCR_DEV_cnt_init[11]), .D (sclear_and_11_dup_158), .CLK (
           CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_7__dup_50 (.Q (FIFO_DEV_count[7]), .D (incdec_mux_7_dup_105)
             , .E (FIFO_DEV_rtlc14_X_0_n123), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_6__dup_51 (.Q (FIFO_DEV_count[6]), .D (incdec_mux_6_dup_104)
             , .E (FIFO_DEV_rtlc14_X_0_n123), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_255_ (.Q (FIFO_DEV_rtlc_msr_n3[255]), .D (
             SIGN_REG_dup_0[7]), .E (nx37353z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_254_ (.Q (FIFO_DEV_rtlc_msr_n3[254]), .D (
             SIGN_REG_dup_0[7]), .E (nx36356z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_253_ (.Q (FIFO_DEV_rtlc_msr_n3[253]), .D (
             SIGN_REG_dup_0[7]), .E (nx35359z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_252_ (.Q (FIFO_DEV_rtlc_msr_n3[252]), .D (
             SIGN_REG_dup_0[7]), .E (nx34362z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_251_ (.Q (FIFO_DEV_rtlc_msr_n3[251]), .D (
             SIGN_REG_dup_0[7]), .E (nx33365z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_250_ (.Q (FIFO_DEV_rtlc_msr_n3[250]), .D (
             SIGN_REG_dup_0[7]), .E (nx32368z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_249_ (.Q (FIFO_DEV_rtlc_msr_n3[249]), .D (
             SIGN_REG_dup_0[7]), .E (nx30372z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_248_ (.Q (FIFO_DEV_rtlc_msr_n3[248]), .D (
             SIGN_REG_dup_0[7]), .E (nx29375z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_247_ (.Q (FIFO_DEV_rtlc_msr_n3[247]), .D (
             SIGN_REG_dup_0[7]), .E (nx28378z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_246_ (.Q (FIFO_DEV_rtlc_msr_n3[246]), .D (
             SIGN_REG_dup_0[7]), .E (nx27381z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_245_ (.Q (FIFO_DEV_rtlc_msr_n3[245]), .D (
             SIGN_REG_dup_0[7]), .E (nx26384z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_244_ (.Q (FIFO_DEV_rtlc_msr_n3[244]), .D (
             SIGN_REG_dup_0[7]), .E (nx25387z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_243_ (.Q (FIFO_DEV_rtlc_msr_n3[243]), .D (
             SIGN_REG_dup_0[7]), .E (nx24390z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_242_ (.Q (FIFO_DEV_rtlc_msr_n3[242]), .D (
             SIGN_REG_dup_0[7]), .E (nx23393z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_241_ (.Q (FIFO_DEV_rtlc_msr_n3[241]), .D (
             SIGN_REG_dup_0[7]), .E (nx22396z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_240_ (.Q (FIFO_DEV_rtlc_msr_n3[240]), .D (
             SIGN_REG_dup_0[7]), .E (nx21399z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_239_ (.Q (FIFO_DEV_rtlc_msr_n3[239]), .D (
             SIGN_REG_dup_0[7]), .E (nx19403z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_238_ (.Q (FIFO_DEV_rtlc_msr_n3[238]), .D (
             SIGN_REG_dup_0[7]), .E (nx18406z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_237_ (.Q (FIFO_DEV_rtlc_msr_n3[237]), .D (
             SIGN_REG_dup_0[7]), .E (nx17409z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_236_ (.Q (FIFO_DEV_rtlc_msr_n3[236]), .D (
             SIGN_REG_dup_0[7]), .E (nx16412z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_235_ (.Q (FIFO_DEV_rtlc_msr_n3[235]), .D (
             SIGN_REG_dup_0[7]), .E (nx15415z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_234_ (.Q (FIFO_DEV_rtlc_msr_n3[234]), .D (
             SIGN_REG_dup_0[7]), .E (nx14418z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_233_ (.Q (FIFO_DEV_rtlc_msr_n3[233]), .D (
             SIGN_REG_dup_0[7]), .E (nx13421z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_232_ (.Q (FIFO_DEV_rtlc_msr_n3[232]), .D (
             SIGN_REG_dup_0[7]), .E (nx12424z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_231_ (.Q (FIFO_DEV_rtlc_msr_n3[231]), .D (
             SIGN_REG_dup_0[7]), .E (nx11427z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_230_ (.Q (FIFO_DEV_rtlc_msr_n3[230]), .D (
             SIGN_REG_dup_0[7]), .E (nx10430z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_229_ (.Q (FIFO_DEV_rtlc_msr_n3[229]), .D (
             SIGN_REG_dup_0[7]), .E (nx8434z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_228_ (.Q (FIFO_DEV_rtlc_msr_n3[228]), .D (
             SIGN_REG_dup_0[7]), .E (nx7437z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_227_ (.Q (FIFO_DEV_rtlc_msr_n3[227]), .D (
             SIGN_REG_dup_0[7]), .E (nx6440z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_226_ (.Q (FIFO_DEV_rtlc_msr_n3[226]), .D (
             SIGN_REG_dup_0[7]), .E (nx5443z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_225_ (.Q (FIFO_DEV_rtlc_msr_n3[225]), .D (
             SIGN_REG_dup_0[7]), .E (nx4446z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_224_ (.Q (FIFO_DEV_rtlc_msr_n3[224]), .D (
             SIGN_REG_dup_0[7]), .E (nx3449z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_223_ (.Q (FIFO_DEV_rtlc_msr_n3[223]), .D (
             SIGN_REG_dup_0[7]), .E (nx2452z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_222_ (.Q (FIFO_DEV_rtlc_msr_n3[222]), .D (
             SIGN_REG_dup_0[7]), .E (nx1455z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_221_ (.Q (FIFO_DEV_rtlc_msr_n3[221]), .D (
             SIGN_REG_dup_0[7]), .E (nx458z1), .CLK (CLK_int), .PRE (RST_int)) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_220_ (.Q (FIFO_DEV_rtlc_msr_n3[220]), .D (
             SIGN_REG_dup_0[7]), .E (nx64997z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_219_ (.Q (FIFO_DEV_rtlc_msr_n3[219]), .D (
             SIGN_REG_dup_0[7]), .E (nx63001z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_218_ (.Q (FIFO_DEV_rtlc_msr_n3[218]), .D (
             SIGN_REG_dup_0[7]), .E (nx62004z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_217_ (.Q (FIFO_DEV_rtlc_msr_n3[217]), .D (
             SIGN_REG_dup_0[7]), .E (nx61007z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_216_ (.Q (FIFO_DEV_rtlc_msr_n3[216]), .D (
             SIGN_REG_dup_0[7]), .E (nx60010z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_215_ (.Q (FIFO_DEV_rtlc_msr_n3[215]), .D (
             SIGN_REG_dup_0[7]), .E (nx59013z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_214_ (.Q (FIFO_DEV_rtlc_msr_n3[214]), .D (
             SIGN_REG_dup_0[7]), .E (nx58016z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_213_ (.Q (FIFO_DEV_rtlc_msr_n3[213]), .D (
             SIGN_REG_dup_0[7]), .E (nx57019z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_212_ (.Q (FIFO_DEV_rtlc_msr_n3[212]), .D (
             SIGN_REG_dup_0[7]), .E (nx56022z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_211_ (.Q (FIFO_DEV_rtlc_msr_n3[211]), .D (
             SIGN_REG_dup_0[7]), .E (nx55025z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_210_ (.Q (FIFO_DEV_rtlc_msr_n3[210]), .D (
             SIGN_REG_dup_0[7]), .E (nx54028z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_209_ (.Q (FIFO_DEV_rtlc_msr_n3[209]), .D (
             SIGN_REG_dup_0[7]), .E (nx52032z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_208_ (.Q (FIFO_DEV_rtlc_msr_n3[208]), .D (
             SIGN_REG_dup_0[7]), .E (nx51035z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_207_ (.Q (FIFO_DEV_rtlc_msr_n3[207]), .D (
             SIGN_REG_dup_0[7]), .E (nx50038z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_206_ (.Q (FIFO_DEV_rtlc_msr_n3[206]), .D (
             SIGN_REG_dup_0[7]), .E (nx49041z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_205_ (.Q (FIFO_DEV_rtlc_msr_n3[205]), .D (
             SIGN_REG_dup_0[7]), .E (nx48044z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_204_ (.Q (FIFO_DEV_rtlc_msr_n3[204]), .D (
             SIGN_REG_dup_0[7]), .E (nx47047z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_203_ (.Q (FIFO_DEV_rtlc_msr_n3[203]), .D (
             SIGN_REG_dup_0[7]), .E (nx46050z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_202_ (.Q (FIFO_DEV_rtlc_msr_n3[202]), .D (
             SIGN_REG_dup_0[7]), .E (nx45053z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_201_ (.Q (FIFO_DEV_rtlc_msr_n3[201]), .D (
             SIGN_REG_dup_0[7]), .E (nx44056z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_200_ (.Q (FIFO_DEV_rtlc_msr_n3[200]), .D (
             SIGN_REG_dup_0[7]), .E (nx43059z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_199_ (.Q (FIFO_DEV_rtlc_msr_n3[199]), .D (
             SIGN_REG_dup_0[7]), .E (nx37436z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_198_ (.Q (FIFO_DEV_rtlc_msr_n3[198]), .D (
             SIGN_REG_dup_0[7]), .E (nx38433z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_197_ (.Q (FIFO_DEV_rtlc_msr_n3[197]), .D (
             SIGN_REG_dup_0[7]), .E (nx39430z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_196_ (.Q (FIFO_DEV_rtlc_msr_n3[196]), .D (
             SIGN_REG_dup_0[7]), .E (nx40427z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_195_ (.Q (FIFO_DEV_rtlc_msr_n3[195]), .D (
             SIGN_REG_dup_0[7]), .E (nx41424z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_194_ (.Q (FIFO_DEV_rtlc_msr_n3[194]), .D (
             SIGN_REG_dup_0[7]), .E (nx42421z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_193_ (.Q (FIFO_DEV_rtlc_msr_n3[193]), .D (
             SIGN_REG_dup_0[7]), .E (nx43418z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_192_ (.Q (FIFO_DEV_rtlc_msr_n3[192]), .D (
             SIGN_REG_dup_0[7]), .E (nx44415z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_191_ (.Q (FIFO_DEV_rtlc_msr_n3[191]), .D (
             SIGN_REG_dup_0[7]), .E (nx45412z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_190_ (.Q (FIFO_DEV_rtlc_msr_n3[190]), .D (
             SIGN_REG_dup_0[7]), .E (nx46409z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_189_ (.Q (FIFO_DEV_rtlc_msr_n3[189]), .D (
             SIGN_REG_dup_0[7]), .E (nx48405z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_188_ (.Q (FIFO_DEV_rtlc_msr_n3[188]), .D (
             SIGN_REG_dup_0[7]), .E (nx49402z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_187_ (.Q (FIFO_DEV_rtlc_msr_n3[187]), .D (
             SIGN_REG_dup_0[7]), .E (nx50399z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_186_ (.Q (FIFO_DEV_rtlc_msr_n3[186]), .D (
             SIGN_REG_dup_0[7]), .E (nx51396z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_185_ (.Q (FIFO_DEV_rtlc_msr_n3[185]), .D (
             SIGN_REG_dup_0[7]), .E (nx52393z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_184_ (.Q (FIFO_DEV_rtlc_msr_n3[184]), .D (
             SIGN_REG_dup_0[7]), .E (nx53390z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_183_ (.Q (FIFO_DEV_rtlc_msr_n3[183]), .D (
             SIGN_REG_dup_0[7]), .E (nx54387z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_182_ (.Q (FIFO_DEV_rtlc_msr_n3[182]), .D (
             SIGN_REG_dup_0[7]), .E (nx55384z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_181_ (.Q (FIFO_DEV_rtlc_msr_n3[181]), .D (
             SIGN_REG_dup_0[7]), .E (nx56381z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_180_ (.Q (FIFO_DEV_rtlc_msr_n3[180]), .D (
             SIGN_REG_dup_0[7]), .E (nx57378z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_179_ (.Q (FIFO_DEV_rtlc_msr_n3[179]), .D (
             SIGN_REG_dup_0[7]), .E (nx59374z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_178_ (.Q (FIFO_DEV_rtlc_msr_n3[178]), .D (
             SIGN_REG_dup_0[7]), .E (nx60371z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_177_ (.Q (FIFO_DEV_rtlc_msr_n3[177]), .D (
             SIGN_REG_dup_0[7]), .E (nx61368z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_176_ (.Q (FIFO_DEV_rtlc_msr_n3[176]), .D (
             SIGN_REG_dup_0[7]), .E (nx62365z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_175_ (.Q (FIFO_DEV_rtlc_msr_n3[175]), .D (
             SIGN_REG_dup_0[7]), .E (nx63362z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_174_ (.Q (FIFO_DEV_rtlc_msr_n3[174]), .D (
             SIGN_REG_dup_0[7]), .E (nx64359z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_173_ (.Q (FIFO_DEV_rtlc_msr_n3[173]), .D (
             SIGN_REG_dup_0[7]), .E (nx65356z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_172_ (.Q (FIFO_DEV_rtlc_msr_n3[172]), .D (
             SIGN_REG_dup_0[7]), .E (nx817z1), .CLK (CLK_int), .PRE (RST_int)) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_171_ (.Q (FIFO_DEV_rtlc_msr_n3[171]), .D (
             SIGN_REG_dup_0[7]), .E (nx1814z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_170_ (.Q (FIFO_DEV_rtlc_msr_n3[170]), .D (
             SIGN_REG_dup_0[7]), .E (nx2811z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_169_ (.Q (FIFO_DEV_rtlc_msr_n3[169]), .D (
             SIGN_REG_dup_0[7]), .E (nx4807z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_168_ (.Q (FIFO_DEV_rtlc_msr_n3[168]), .D (
             SIGN_REG_dup_0[7]), .E (nx5804z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_167_ (.Q (FIFO_DEV_rtlc_msr_n3[167]), .D (
             SIGN_REG_dup_0[7]), .E (nx6801z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_166_ (.Q (FIFO_DEV_rtlc_msr_n3[166]), .D (
             SIGN_REG_dup_0[7]), .E (nx7798z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_165_ (.Q (FIFO_DEV_rtlc_msr_n3[165]), .D (
             SIGN_REG_dup_0[7]), .E (nx8795z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_164_ (.Q (FIFO_DEV_rtlc_msr_n3[164]), .D (
             SIGN_REG_dup_0[7]), .E (nx9792z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_163_ (.Q (FIFO_DEV_rtlc_msr_n3[163]), .D (
             SIGN_REG_dup_0[7]), .E (nx10789z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_162_ (.Q (FIFO_DEV_rtlc_msr_n3[162]), .D (
             SIGN_REG_dup_0[7]), .E (nx11786z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_161_ (.Q (FIFO_DEV_rtlc_msr_n3[161]), .D (
             SIGN_REG_dup_0[7]), .E (nx12783z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_160_ (.Q (FIFO_DEV_rtlc_msr_n3[160]), .D (
             SIGN_REG_dup_0[7]), .E (nx13780z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_159_ (.Q (FIFO_DEV_rtlc_msr_n3[159]), .D (
             SIGN_REG_dup_0[7]), .E (nx15776z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_158_ (.Q (FIFO_DEV_rtlc_msr_n3[158]), .D (
             SIGN_REG_dup_0[7]), .E (nx16773z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_157_ (.Q (FIFO_DEV_rtlc_msr_n3[157]), .D (
             SIGN_REG_dup_0[7]), .E (nx17770z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_156_ (.Q (FIFO_DEV_rtlc_msr_n3[156]), .D (
             SIGN_REG_dup_0[7]), .E (nx18767z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_155_ (.Q (FIFO_DEV_rtlc_msr_n3[155]), .D (
             SIGN_REG_dup_0[7]), .E (nx19764z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_154_ (.Q (FIFO_DEV_rtlc_msr_n3[154]), .D (
             SIGN_REG_dup_0[7]), .E (nx20761z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_153_ (.Q (FIFO_DEV_rtlc_msr_n3[153]), .D (
             SIGN_REG_dup_0[7]), .E (nx21758z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_152_ (.Q (FIFO_DEV_rtlc_msr_n3[152]), .D (
             SIGN_REG_dup_0[7]), .E (nx22755z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_151_ (.Q (FIFO_DEV_rtlc_msr_n3[151]), .D (
             SIGN_REG_dup_0[7]), .E (nx23752z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_150_ (.Q (FIFO_DEV_rtlc_msr_n3[150]), .D (
             SIGN_REG_dup_0[7]), .E (nx24749z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_149_ (.Q (FIFO_DEV_rtlc_msr_n3[149]), .D (
             SIGN_REG_dup_0[7]), .E (nx26745z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_148_ (.Q (FIFO_DEV_rtlc_msr_n3[148]), .D (
             SIGN_REG_dup_0[7]), .E (nx27742z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_147_ (.Q (FIFO_DEV_rtlc_msr_n3[147]), .D (
             SIGN_REG_dup_0[7]), .E (nx28739z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_146_ (.Q (FIFO_DEV_rtlc_msr_n3[146]), .D (
             SIGN_REG_dup_0[7]), .E (nx29736z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_145_ (.Q (FIFO_DEV_rtlc_msr_n3[145]), .D (
             SIGN_REG_dup_0[7]), .E (nx30733z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_144_ (.Q (FIFO_DEV_rtlc_msr_n3[144]), .D (
             SIGN_REG_dup_0[7]), .E (nx31730z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_143_ (.Q (FIFO_DEV_rtlc_msr_n3[143]), .D (
             SIGN_REG_dup_0[7]), .E (nx32727z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_142_ (.Q (FIFO_DEV_rtlc_msr_n3[142]), .D (
             SIGN_REG_dup_0[7]), .E (nx33724z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_141_ (.Q (FIFO_DEV_rtlc_msr_n3[141]), .D (
             SIGN_REG_dup_0[7]), .E (nx34721z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_140_ (.Q (FIFO_DEV_rtlc_msr_n3[140]), .D (
             SIGN_REG_dup_0[7]), .E (nx35718z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_139_ (.Q (FIFO_DEV_rtlc_msr_n3[139]), .D (
             SIGN_REG_dup_0[7]), .E (nx37714z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_138_ (.Q (FIFO_DEV_rtlc_msr_n3[138]), .D (
             SIGN_REG_dup_0[7]), .E (nx38711z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_137_ (.Q (FIFO_DEV_rtlc_msr_n3[137]), .D (
             SIGN_REG_dup_0[7]), .E (nx39708z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_136_ (.Q (FIFO_DEV_rtlc_msr_n3[136]), .D (
             SIGN_REG_dup_0[7]), .E (nx40705z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_135_ (.Q (FIFO_DEV_rtlc_msr_n3[135]), .D (
             SIGN_REG_dup_0[7]), .E (nx41702z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_134_ (.Q (FIFO_DEV_rtlc_msr_n3[134]), .D (
             SIGN_REG_dup_0[7]), .E (nx42699z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_133_ (.Q (FIFO_DEV_rtlc_msr_n3[133]), .D (
             SIGN_REG_dup_0[7]), .E (nx43696z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_132_ (.Q (FIFO_DEV_rtlc_msr_n3[132]), .D (
             SIGN_REG_dup_0[7]), .E (nx44693z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_131_ (.Q (FIFO_DEV_rtlc_msr_n3[131]), .D (
             SIGN_REG_dup_0[7]), .E (nx45690z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_130_ (.Q (FIFO_DEV_rtlc_msr_n3[130]), .D (
             SIGN_REG_dup_0[7]), .E (nx46687z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_129_ (.Q (FIFO_DEV_rtlc_msr_n3[129]), .D (
             SIGN_REG_dup_0[7]), .E (nx48683z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_128_ (.Q (FIFO_DEV_rtlc_msr_n3[128]), .D (
             SIGN_REG_dup_0[7]), .E (nx49680z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_127_ (.Q (FIFO_DEV_rtlc_msr_n3[127]), .D (
             SIGN_REG_dup_0[7]), .E (nx50677z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_126_ (.Q (FIFO_DEV_rtlc_msr_n3[126]), .D (
             SIGN_REG_dup_0[7]), .E (nx51674z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_125_ (.Q (FIFO_DEV_rtlc_msr_n3[125]), .D (
             SIGN_REG_dup_0[7]), .E (nx52671z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_124_ (.Q (FIFO_DEV_rtlc_msr_n3[124]), .D (
             SIGN_REG_dup_0[7]), .E (nx53668z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_123_ (.Q (FIFO_DEV_rtlc_msr_n3[123]), .D (
             SIGN_REG_dup_0[7]), .E (nx54665z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_122_ (.Q (FIFO_DEV_rtlc_msr_n3[122]), .D (
             SIGN_REG_dup_0[7]), .E (nx55662z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_121_ (.Q (FIFO_DEV_rtlc_msr_n3[121]), .D (
             SIGN_REG_dup_0[7]), .E (nx56659z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_120_ (.Q (FIFO_DEV_rtlc_msr_n3[120]), .D (
             SIGN_REG_dup_0[7]), .E (nx57656z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_119_ (.Q (FIFO_DEV_rtlc_msr_n3[119]), .D (
             SIGN_REG_dup_0[7]), .E (nx59652z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_118_ (.Q (FIFO_DEV_rtlc_msr_n3[118]), .D (
             SIGN_REG_dup_0[7]), .E (nx60649z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_117_ (.Q (FIFO_DEV_rtlc_msr_n3[117]), .D (
             SIGN_REG_dup_0[7]), .E (nx61646z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_116_ (.Q (FIFO_DEV_rtlc_msr_n3[116]), .D (
             SIGN_REG_dup_0[7]), .E (nx62643z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_115_ (.Q (FIFO_DEV_rtlc_msr_n3[115]), .D (
             SIGN_REG_dup_0[7]), .E (nx63640z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_114_ (.Q (FIFO_DEV_rtlc_msr_n3[114]), .D (
             SIGN_REG_dup_0[7]), .E (nx64637z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_113_ (.Q (FIFO_DEV_rtlc_msr_n3[113]), .D (
             SIGN_REG_dup_0[7]), .E (nx98z1), .CLK (CLK_int), .PRE (RST_int)) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_112_ (.Q (FIFO_DEV_rtlc_msr_n3[112]), .D (
             SIGN_REG_dup_0[7]), .E (nx1095z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_111_ (.Q (FIFO_DEV_rtlc_msr_n3[111]), .D (
             SIGN_REG_dup_0[7]), .E (nx2092z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_110_ (.Q (FIFO_DEV_rtlc_msr_n3[110]), .D (
             SIGN_REG_dup_0[7]), .E (nx3089z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_109_ (.Q (FIFO_DEV_rtlc_msr_n3[109]), .D (
             SIGN_REG_dup_0[7]), .E (nx5085z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_108_ (.Q (FIFO_DEV_rtlc_msr_n3[108]), .D (
             SIGN_REG_dup_0[7]), .E (nx6082z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_107_ (.Q (FIFO_DEV_rtlc_msr_n3[107]), .D (
             SIGN_REG_dup_0[7]), .E (nx7079z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_106_ (.Q (FIFO_DEV_rtlc_msr_n3[106]), .D (
             SIGN_REG_dup_0[7]), .E (nx8076z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_105_ (.Q (FIFO_DEV_rtlc_msr_n3[105]), .D (
             SIGN_REG_dup_0[7]), .E (nx9073z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_104_ (.Q (FIFO_DEV_rtlc_msr_n3[104]), .D (
             SIGN_REG_dup_0[7]), .E (nx10070z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_103_ (.Q (FIFO_DEV_rtlc_msr_n3[103]), .D (
             SIGN_REG_dup_0[7]), .E (nx11067z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_102_ (.Q (FIFO_DEV_rtlc_msr_n3[102]), .D (
             SIGN_REG_dup_0[7]), .E (nx12064z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_101_ (.Q (FIFO_DEV_rtlc_msr_n3[101]), .D (
             SIGN_REG_dup_0[7]), .E (nx13061z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_100_ (.Q (FIFO_DEV_rtlc_msr_n3[100]), .D (
             SIGN_REG_dup_0[7]), .E (nx14058z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_99_ (.Q (FIFO_DEV_rtlc_msr_n3[99]), .D (
             SIGN_REG_dup_0[7]), .E (nx5577z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_98_ (.Q (FIFO_DEV_rtlc_msr_n3[98]), .D (
             SIGN_REG_dup_0[7]), .E (nx6574z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_97_ (.Q (FIFO_DEV_rtlc_msr_n3[97]), .D (
             SIGN_REG_dup_0[7]), .E (nx7571z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_96_ (.Q (FIFO_DEV_rtlc_msr_n3[96]), .D (
             SIGN_REG_dup_0[7]), .E (nx8568z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_95_ (.Q (FIFO_DEV_rtlc_msr_n3[95]), .D (
             SIGN_REG_dup_0[7]), .E (nx9565z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_94_ (.Q (FIFO_DEV_rtlc_msr_n3[94]), .D (
             SIGN_REG_dup_0[7]), .E (nx10562z4), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_93_ (.Q (FIFO_DEV_rtlc_msr_n3[93]), .D (
             SIGN_REG_dup_0[7]), .E (nx11559z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_92_ (.Q (FIFO_DEV_rtlc_msr_n3[92]), .D (
             SIGN_REG_dup_0[7]), .E (nx12556z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_91_ (.Q (FIFO_DEV_rtlc_msr_n3[91]), .D (
             SIGN_REG_dup_0[7]), .E (nx13553z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_90_ (.Q (FIFO_DEV_rtlc_msr_n3[90]), .D (
             SIGN_REG_dup_0[7]), .E (nx14550z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_89_ (.Q (FIFO_DEV_rtlc_msr_n3[89]), .D (
             SIGN_REG_dup_0[7]), .E (nx16546z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_88_ (.Q (FIFO_DEV_rtlc_msr_n3[88]), .D (
             SIGN_REG_dup_0[7]), .E (nx17543z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_87_ (.Q (FIFO_DEV_rtlc_msr_n3[87]), .D (
             SIGN_REG_dup_0[7]), .E (nx18540z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_86_ (.Q (FIFO_DEV_rtlc_msr_n3[86]), .D (
             SIGN_REG_dup_0[7]), .E (nx19537z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_85_ (.Q (FIFO_DEV_rtlc_msr_n3[85]), .D (
             SIGN_REG_dup_0[7]), .E (nx20534z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_84_ (.Q (FIFO_DEV_rtlc_msr_n3[84]), .D (
             SIGN_REG_dup_0[7]), .E (nx21531z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_83_ (.Q (FIFO_DEV_rtlc_msr_n3[83]), .D (
             SIGN_REG_dup_0[7]), .E (nx22528z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_82_ (.Q (FIFO_DEV_rtlc_msr_n3[82]), .D (
             SIGN_REG_dup_0[7]), .E (nx23525z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_81_ (.Q (FIFO_DEV_rtlc_msr_n3[81]), .D (
             SIGN_REG_dup_0[7]), .E (nx24522z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_80_ (.Q (FIFO_DEV_rtlc_msr_n3[80]), .D (
             SIGN_REG_dup_0[7]), .E (nx25519z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_79_ (.Q (FIFO_DEV_rtlc_msr_n3[79]), .D (
             SIGN_REG_dup_0[7]), .E (nx27515z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_78_ (.Q (FIFO_DEV_rtlc_msr_n3[78]), .D (
             SIGN_REG_dup_0[7]), .E (nx28512z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_77_ (.Q (FIFO_DEV_rtlc_msr_n3[77]), .D (
             SIGN_REG_dup_0[7]), .E (nx29509z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_76_ (.Q (FIFO_DEV_rtlc_msr_n3[76]), .D (
             SIGN_REG_dup_0[7]), .E (nx30506z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_75_ (.Q (FIFO_DEV_rtlc_msr_n3[75]), .D (
             SIGN_REG_dup_0[7]), .E (nx31503z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_74_ (.Q (FIFO_DEV_rtlc_msr_n3[74]), .D (
             SIGN_REG_dup_0[7]), .E (nx32500z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_73_ (.Q (FIFO_DEV_rtlc_msr_n3[73]), .D (
             SIGN_REG_dup_0[7]), .E (nx33497z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_72_ (.Q (FIFO_DEV_rtlc_msr_n3[72]), .D (
             SIGN_REG_dup_0[7]), .E (nx34494z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_71_ (.Q (FIFO_DEV_rtlc_msr_n3[71]), .D (
             SIGN_REG_dup_0[7]), .E (nx35491z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_70_ (.Q (FIFO_DEV_rtlc_msr_n3[70]), .D (
             SIGN_REG_dup_0[7]), .E (nx36488z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_69_ (.Q (FIFO_DEV_rtlc_msr_n3[69]), .D (
             SIGN_REG_dup_0[7]), .E (nx38484z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_68_ (.Q (FIFO_DEV_rtlc_msr_n3[68]), .D (
             SIGN_REG_dup_0[7]), .E (nx39481z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_67_ (.Q (FIFO_DEV_rtlc_msr_n3[67]), .D (
             SIGN_REG_dup_0[7]), .E (nx40478z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_66_ (.Q (FIFO_DEV_rtlc_msr_n3[66]), .D (
             SIGN_REG_dup_0[7]), .E (nx41475z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_65_ (.Q (FIFO_DEV_rtlc_msr_n3[65]), .D (
             SIGN_REG_dup_0[7]), .E (nx42472z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_64_ (.Q (FIFO_DEV_rtlc_msr_n3[64]), .D (
             SIGN_REG_dup_0[7]), .E (nx43469z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_63_ (.Q (FIFO_DEV_rtlc_msr_n3[63]), .D (
             SIGN_REG_dup_0[7]), .E (nx44466z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_62_ (.Q (FIFO_DEV_rtlc_msr_n3[62]), .D (
             SIGN_REG_dup_0[7]), .E (nx45463z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_61_ (.Q (FIFO_DEV_rtlc_msr_n3[61]), .D (
             SIGN_REG_dup_0[7]), .E (nx46460z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_60_ (.Q (FIFO_DEV_rtlc_msr_n3[60]), .D (
             SIGN_REG_dup_0[7]), .E (nx47457z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_59_ (.Q (FIFO_DEV_rtlc_msr_n3[59]), .D (
             SIGN_REG_dup_0[7]), .E (nx49453z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_58_ (.Q (FIFO_DEV_rtlc_msr_n3[58]), .D (
             SIGN_REG_dup_0[7]), .E (nx50450z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_57_ (.Q (FIFO_DEV_rtlc_msr_n3[57]), .D (
             SIGN_REG_dup_0[7]), .E (nx51447z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_56_ (.Q (FIFO_DEV_rtlc_msr_n3[56]), .D (
             SIGN_REG_dup_0[7]), .E (nx52444z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_55_ (.Q (FIFO_DEV_rtlc_msr_n3[55]), .D (
             SIGN_REG_dup_0[7]), .E (nx53441z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_54_ (.Q (FIFO_DEV_rtlc_msr_n3[54]), .D (
             SIGN_REG_dup_0[7]), .E (nx54438z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_53_ (.Q (FIFO_DEV_rtlc_msr_n3[53]), .D (
             SIGN_REG_dup_0[7]), .E (nx55435z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_52_ (.Q (FIFO_DEV_rtlc_msr_n3[52]), .D (
             SIGN_REG_dup_0[7]), .E (nx56432z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_51_ (.Q (FIFO_DEV_rtlc_msr_n3[51]), .D (
             SIGN_REG_dup_0[7]), .E (nx57429z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_50_ (.Q (FIFO_DEV_rtlc_msr_n3[50]), .D (
             SIGN_REG_dup_0[7]), .E (nx58426z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_49_ (.Q (FIFO_DEV_rtlc_msr_n3[49]), .D (
             SIGN_REG_dup_0[7]), .E (nx60422z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_48_ (.Q (FIFO_DEV_rtlc_msr_n3[48]), .D (
             SIGN_REG_dup_0[7]), .E (nx61419z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_47_ (.Q (FIFO_DEV_rtlc_msr_n3[47]), .D (
             SIGN_REG_dup_0[7]), .E (nx62416z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_46_ (.Q (FIFO_DEV_rtlc_msr_n3[46]), .D (
             SIGN_REG_dup_0[7]), .E (nx63413z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_45_ (.Q (FIFO_DEV_rtlc_msr_n3[45]), .D (
             SIGN_REG_dup_0[7]), .E (nx64410z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_44_ (.Q (FIFO_DEV_rtlc_msr_n3[44]), .D (
             SIGN_REG_dup_0[7]), .E (nx65407z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_43_ (.Q (FIFO_DEV_rtlc_msr_n3[43]), .D (
             SIGN_REG_dup_0[7]), .E (nx868z1), .CLK (CLK_int), .PRE (RST_int)) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_42_ (.Q (FIFO_DEV_rtlc_msr_n3[42]), .D (
             SIGN_REG_dup_0[7]), .E (nx1865z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_41_ (.Q (FIFO_DEV_rtlc_msr_n3[41]), .D (
             SIGN_REG_dup_0[7]), .E (nx2862z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_40_ (.Q (FIFO_DEV_rtlc_msr_n3[40]), .D (
             SIGN_REG_dup_0[7]), .E (nx3859z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_39_ (.Q (FIFO_DEV_rtlc_msr_n3[39]), .D (
             SIGN_REG_dup_0[7]), .E (nx5855z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_38_ (.Q (FIFO_DEV_rtlc_msr_n3[38]), .D (
             SIGN_REG_dup_0[7]), .E (nx6852z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_37_ (.Q (FIFO_DEV_rtlc_msr_n3[37]), .D (
             SIGN_REG_dup_0[7]), .E (nx7849z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_36_ (.Q (FIFO_DEV_rtlc_msr_n3[36]), .D (
             SIGN_REG_dup_0[7]), .E (nx8846z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_35_ (.Q (FIFO_DEV_rtlc_msr_n3[35]), .D (
             SIGN_REG_dup_0[7]), .E (nx9843z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_34_ (.Q (FIFO_DEV_rtlc_msr_n3[34]), .D (
             SIGN_REG_dup_0[7]), .E (nx10840z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_33_ (.Q (FIFO_DEV_rtlc_msr_n3[33]), .D (
             SIGN_REG_dup_0[7]), .E (nx11837z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_32_ (.Q (FIFO_DEV_rtlc_msr_n3[32]), .D (
             SIGN_REG_dup_0[7]), .E (nx12834z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_31_ (.Q (FIFO_DEV_rtlc_msr_n3[31]), .D (
             SIGN_REG_dup_0[7]), .E (nx13831z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_30_ (.Q (FIFO_DEV_rtlc_msr_n3[30]), .D (
             SIGN_REG_dup_0[7]), .E (nx14828z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_29_ (.Q (FIFO_DEV_rtlc_msr_n3[29]), .D (
             SIGN_REG_dup_0[7]), .E (nx16824z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_28_ (.Q (FIFO_DEV_rtlc_msr_n3[28]), .D (
             SIGN_REG_dup_0[7]), .E (nx17821z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_27_ (.Q (FIFO_DEV_rtlc_msr_n3[27]), .D (
             SIGN_REG_dup_0[7]), .E (nx18818z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_26_ (.Q (FIFO_DEV_rtlc_msr_n3[26]), .D (
             SIGN_REG_dup_0[7]), .E (nx19815z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_25_ (.Q (FIFO_DEV_rtlc_msr_n3[25]), .D (
             SIGN_REG_dup_0[7]), .E (nx20812z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_24_ (.Q (FIFO_DEV_rtlc_msr_n3[24]), .D (
             SIGN_REG_dup_0[7]), .E (nx21809z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_23_ (.Q (FIFO_DEV_rtlc_msr_n3[23]), .D (
             SIGN_REG_dup_0[7]), .E (nx22806z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_22_ (.Q (FIFO_DEV_rtlc_msr_n3[22]), .D (
             SIGN_REG_dup_0[7]), .E (nx23803z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_21_ (.Q (FIFO_DEV_rtlc_msr_n3[21]), .D (
             SIGN_REG_dup_0[7]), .E (nx24800z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_20_ (.Q (FIFO_DEV_rtlc_msr_n3[20]), .D (
             SIGN_REG_dup_0[7]), .E (nx25797z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_19_ (.Q (FIFO_DEV_rtlc_msr_n3[19]), .D (
             SIGN_REG_dup_0[7]), .E (nx27793z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_18_ (.Q (FIFO_DEV_rtlc_msr_n3[18]), .D (
             SIGN_REG_dup_0[7]), .E (nx28790z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_17_ (.Q (FIFO_DEV_rtlc_msr_n3[17]), .D (
             SIGN_REG_dup_0[7]), .E (nx29787z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_16_ (.Q (FIFO_DEV_rtlc_msr_n3[16]), .D (
             SIGN_REG_dup_0[7]), .E (nx30784z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_15_ (.Q (FIFO_DEV_rtlc_msr_n3[15]), .D (
             SIGN_REG_dup_0[7]), .E (nx31781z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_14_ (.Q (FIFO_DEV_rtlc_msr_n3[14]), .D (
             SIGN_REG_dup_0[7]), .E (nx32778z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_13_ (.Q (FIFO_DEV_rtlc_msr_n3[13]), .D (
             SIGN_REG_dup_0[7]), .E (nx33775z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_12_ (.Q (FIFO_DEV_rtlc_msr_n3[12]), .D (
             SIGN_REG_dup_0[7]), .E (nx34772z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_11_ (.Q (FIFO_DEV_rtlc_msr_n3[11]), .D (
             SIGN_REG_dup_0[7]), .E (nx35769z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_10_ (.Q (FIFO_DEV_rtlc_msr_n3[10]), .D (
             SIGN_REG_dup_0[7]), .E (nx36766z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_9_ (.Q (FIFO_DEV_rtlc_msr_n3[9]), .D (
             SIGN_REG_dup_0[7]), .E (nx48358z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_8_ (.Q (FIFO_DEV_rtlc_msr_n3[8]), .D (
             SIGN_REG_dup_0[7]), .E (nx47361z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_7_ (.Q (FIFO_DEV_rtlc_msr_n3[7]), .D (
             SIGN_REG_dup_0[7]), .E (nx46364z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_6_ (.Q (FIFO_DEV_rtlc_msr_n3[6]), .D (
             SIGN_REG_dup_0[7]), .E (nx45367z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_5_ (.Q (FIFO_DEV_rtlc_msr_n3[5]), .D (
             SIGN_REG_dup_0[7]), .E (nx44370z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_4_ (.Q (FIFO_DEV_rtlc_msr_n3[4]), .D (
             SIGN_REG_dup_0[7]), .E (nx43373z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_3_ (.Q (FIFO_DEV_rtlc_msr_n3[3]), .D (
             SIGN_REG_dup_0[7]), .E (nx42376z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_2_ (.Q (FIFO_DEV_rtlc_msr_n3[2]), .D (
             SIGN_REG_dup_0[7]), .E (nx41379z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_1_ (.Q (FIFO_DEV_rtlc_msr_n3[1]), .D (
             SIGN_REG_dup_0[7]), .E (nx40382z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1E0P0 FIFO_DEV_reg_rtlc_msr_n3_0_ (.Q (FIFO_DEV_rtlc_msr_n3[0]), .D (
             SIGN_REG_dup_0[7]), .E (nx39385z1), .CLK (CLK_int), .PRE (RST_int)
             ) ;
    DFN1C0 ENCR_DEV_reg_strob_data_tmp (.Q (ENCR_DEV_strob_data_tmp), .D (
           STB_DATA_int), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1P0 ENCR_DEV_reg_prev_0_ (.Q (ENCR_DEV_prev[0]), .D (nx7516z1), .CLK (
           CLK_int), .PRE (RST_int)) ;
    DFN1E0C0 ENCR_DEV_modgen_counter_key_cnt_reg_q_1_ (.Q (ENCR_DEV_key_cnt[1])
             , .D (nx44635z1), .E (nx45632z2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_modgen_counter_key_cnt_reg_q_0_ (.Q (ENCR_DEV_key_cnt[0])
             , .D (nx45632z1), .E (nx45632z2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_prev_7_ (.Q (ENCR_DEV_prev[7]), .D (nx14495z1), .CLK (
           CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_19_ (.Q (ENCR_DEV_err_cnt[19]), .D (sclear_and_19_dup_738), .E (
             nx25368z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_18_ (.Q (ENCR_DEV_err_cnt[18]), .D (sclear_and_18_dup_737), .E (
             nx25368z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_23_ (.Q (ENCR_DEV_err_cnt[23]), .D (sclear_and_23_dup_742), .E (
             nx25368z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_22_ (.Q (ENCR_DEV_err_cnt[22]), .D (sclear_and_22_dup_741), .E (
             nx25368z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_5__dup_6 (.Q (ENCR_DEV_err_cnt[5]), .D (sclear_and_5_dup_724)
             , .E (nx25368z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_4__dup_7 (.Q (ENCR_DEV_err_cnt[4]), .D (sclear_and_4_dup_723)
             , .E (nx25368z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_7__dup_4 (.Q (ENCR_DEV_err_cnt[7]), .D (sclear_and_7_dup_726)
             , .E (nx25368z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_6__dup_5 (.Q (ENCR_DEV_err_cnt[6]), .D (sclear_and_6_dup_725)
             , .E (nx25368z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_3__dup_8 (.Q (ENCR_DEV_err_cnt[3]), .D (sclear_and_3_dup_722)
             , .E (nx25368z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_2__dup_9 (.Q (ENCR_DEV_err_cnt[2]), .D (sclear_and_2_dup_721)
             , .E (nx25368z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_1__dup_10 (.Q (ENCR_DEV_err_cnt[1]), .D (sclear_and_1_dup_720
             ), .E (nx25368z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_63_ (.Q (ENCR_DEV_err_cnt[63]), .D (sclear_and_63_dup_782), .E (
             nx25368z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_61_ (.Q (ENCR_DEV_err_cnt[61]), .D (sclear_and_61_dup_780), .E (
             nx25368z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_62_ (.Q (ENCR_DEV_err_cnt[62]), .D (sclear_and_62_dup_781), .E (
             ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_4__dup_28 (.Q (ENCR_DEV_encry_cnt[4]), .D (
             sclear_and_4_dup_118), .E (ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int
             ), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_3__dup_29 (.Q (ENCR_DEV_encry_cnt[3]), .D (
             sclear_and_3_dup_117), .E (ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int
             ), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_8__dup_24 (.Q (ENCR_DEV_encry_cnt[8]), .D (
             sclear_and_8_dup_122), .E (ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int
             ), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_7__dup_25 (.Q (ENCR_DEV_encry_cnt[7]), .D (
             sclear_and_7_dup_121), .E (ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int
             ), .CLR (RST_int)) ;
    DFN1C0 reg_q_10_ (.Q (ENCR_DEV_cnt_init[10]), .D (sclear_and_10_dup_157), .CLK (
           CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_58_ (.Q (ENCR_DEV_reg_str_1[58]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[58]), .E (nx19668z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1C0 ENCR_DEV_reg_data_reg_7_ (.Q (ENCR_DEV_data_reg[7]), .D (DATA_int[7])
           , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_103_ (.Q (ENCR_DEV_reg_str_3[103]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[103]), .E (nx55223z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_85_ (.Q (ENCR_DEV_reg_str_1[85]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[85]), .E (nx55223z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_76_ (.Q (ENCR_DEV_reg_str_2[76]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[76]), .E (nx19668z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_59_ (.Q (ENCR_DEV_reg_str_1[59]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[59]), .E (nx19668z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1C0 ENCR_DEV_reg_data_reg_6_ (.Q (ENCR_DEV_data_reg[6]), .D (DATA_int[6])
           , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_59_ (.Q (ENCR_DEV_reg_str_3[59]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[59]), .E (nx55223z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_86_ (.Q (ENCR_DEV_reg_str_1[86]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[86]), .E (nx55223z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_77_ (.Q (ENCR_DEV_reg_str_2[77]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[77]), .E (nx19668z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_60_ (.Q (ENCR_DEV_reg_str_1[60]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[60]), .E (nx19668z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1C0 ENCR_DEV_reg_data_reg_5_ (.Q (ENCR_DEV_data_reg[5]), .D (DATA_int[5])
           , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_105_ (.Q (ENCR_DEV_reg_str_3[105]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[105]), .E (nx55223z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_87_ (.Q (ENCR_DEV_reg_str_1[87]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[87]), .E (nx55223z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_78_ (.Q (ENCR_DEV_reg_str_2[78]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[78]), .E (nx19668z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_61_ (.Q (ENCR_DEV_reg_str_1[61]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[61]), .E (nx19668z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1C0 ENCR_DEV_reg_data_reg_4_ (.Q (ENCR_DEV_data_reg[4]), .D (DATA_int[4])
           , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_88_ (.Q (ENCR_DEV_reg_str_1[88]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[88]), .E (nx55223z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_79_ (.Q (ENCR_DEV_reg_str_2[79]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[79]), .E (nx19668z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_106_ (.Q (ENCR_DEV_reg_str_3[106]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[106]), .E (
             NOT_ENCR_DEV_rtlc15n968__repl4), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_62_ (.Q (ENCR_DEV_reg_str_1[62]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[62]), .E (nx19668z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1C0 ENCR_DEV_reg_data_reg_3_ (.Q (ENCR_DEV_data_reg[3]), .D (DATA_int[3])
           , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_89_ (.Q (ENCR_DEV_reg_str_1[89]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[89]), .E (NOT_ENCR_DEV_rtlc15n968__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_80_ (.Q (ENCR_DEV_reg_str_2[80]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[80]), .E (NOT_ENCR_DEV_rtlc15n968__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_107_ (.Q (ENCR_DEV_reg_str_3[107]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[107]), .E (
             NOT_ENCR_DEV_rtlc15n968__repl4), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_63_ (.Q (ENCR_DEV_reg_str_1[63]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[63]), .E (nx19668z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1C0 ENCR_DEV_reg_data_reg_2_ (.Q (ENCR_DEV_data_reg[2]), .D (DATA_int[2])
           , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_108_ (.Q (ENCR_DEV_reg_str_3[108]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[108]), .E (nx19668z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_90_ (.Q (ENCR_DEV_reg_str_1[90]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[90]), .E (NOT_ENCR_DEV_rtlc15n968__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_81_ (.Q (ENCR_DEV_reg_str_2[81]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[81]), .E (NOT_ENCR_DEV_rtlc15n968__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_64_ (.Q (ENCR_DEV_reg_str_1[64]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[64]), .E (nx19668z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1C0 ENCR_DEV_reg_data_reg_1_ (.Q (ENCR_DEV_data_reg[1]), .D (DATA_int[1])
           , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_109_ (.Q (ENCR_DEV_reg_str_3[109]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[109]), .E (nx19668z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_91_ (.Q (ENCR_DEV_reg_str_1[91]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[91]), .E (NOT_ENCR_DEV_rtlc15n968__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_82_ (.Q (ENCR_DEV_reg_str_2[82]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[82]), .E (NOT_ENCR_DEV_rtlc15n968__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_68_ (.Q (ENCR_DEV_reg_str_2[68]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[68]), .E (nx19668z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1C0 ENCR_DEV_reg_data_reg_0_ (.Q (ENCR_DEV_data_reg[0]), .D (DATA_int[0])
           , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_65_ (.Q (ENCR_DEV_reg_str_3[65]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[65]), .E (NOT_ENCR_DEV_rtlc15n968__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_65_ (.Q (ENCR_DEV_reg_str_1[65]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[65]), .E (nx19668z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_83_ (.Q (ENCR_DEV_reg_str_2[83]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[83]), .E (NOT_ENCR_DEV_rtlc15n968__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_27_ (.Q (ENCR_DEV_err_cnt[27]), .D (sclear_and_27_dup_746), .E (
             ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_26_ (.Q (ENCR_DEV_err_cnt[26]), .D (sclear_and_26_dup_745), .E (
             ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_31_ (.Q (ENCR_DEV_err_cnt[31]), .D (sclear_and_31_dup_750), .E (
             ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_30_ (.Q (ENCR_DEV_err_cnt[30]), .D (sclear_and_30_dup_749), .E (
             ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_17_ (.Q (ENCR_DEV_err_cnt[17]), .D (sclear_and_17_dup_736), .E (
             ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_16_ (.Q (ENCR_DEV_err_cnt[16]), .D (sclear_and_16_dup_735), .E (
             ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_21_ (.Q (ENCR_DEV_err_cnt[21]), .D (sclear_and_21_dup_740), .E (
             ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_20_ (.Q (ENCR_DEV_err_cnt[20]), .D (sclear_and_20_dup_739), .E (
             ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_35_ (.Q (ENCR_DEV_err_cnt[35]), .D (sclear_and_35_dup_754), .E (
             ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_34_ (.Q (ENCR_DEV_err_cnt[34]), .D (sclear_and_34_dup_753), .E (
             ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_39_ (.Q (ENCR_DEV_err_cnt[39]), .D (sclear_and_39_dup_758), .E (
             ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_38_ (.Q (ENCR_DEV_err_cnt[38]), .D (sclear_and_38_dup_757), .E (
             ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_43_ (.Q (ENCR_DEV_err_cnt[43]), .D (sclear_and_43_dup_762), .E (
             ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_42_ (.Q (ENCR_DEV_err_cnt[42]), .D (sclear_and_42_dup_761), .E (
             ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_47_ (.Q (ENCR_DEV_err_cnt[47]), .D (sclear_and_47_dup_766), .E (
             ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_46_ (.Q (ENCR_DEV_err_cnt[46]), .D (sclear_and_46_dup_765), .E (
             ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_11__dup_0 (.Q (ENCR_DEV_err_cnt[11]), .D (
             sclear_and_11_dup_730), .E (ENCR_DEV_rtlcn483__repl2), .CLK (
             CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_10__dup_1 (.Q (ENCR_DEV_err_cnt[10]), .D (
             sclear_and_10_dup_729), .E (ENCR_DEV_rtlcn483__repl2), .CLK (
             CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_15_ (.Q (ENCR_DEV_err_cnt[15]), .D (sclear_and_15_dup_734), .E (
             ENCR_DEV_rtlcn483__repl2), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_14_ (.Q (ENCR_DEV_err_cnt[14]), .D (sclear_and_14_dup_733), .E (
             ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_60_ (.Q (ENCR_DEV_err_cnt[60]), .D (sclear_and_60_dup_779), .E (
             ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_0__dup_11 (.Q (ENCR_DEV_err_cnt[0]), .D (sclear_and_0_dup_719
             ), .E (ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_51_ (.Q (ENCR_DEV_err_cnt[51]), .D (sclear_and_51_dup_770), .E (
             ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_50_ (.Q (ENCR_DEV_err_cnt[50]), .D (sclear_and_50_dup_769), .E (
             ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_55_ (.Q (ENCR_DEV_err_cnt[55]), .D (sclear_and_55_dup_774), .E (
             ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_54_ (.Q (ENCR_DEV_err_cnt[54]), .D (sclear_and_54_dup_773), .E (
             ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_59_ (.Q (ENCR_DEV_err_cnt[59]), .D (sclear_and_59_dup_778), .E (
             ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_58_ (.Q (ENCR_DEV_err_cnt[58]), .D (sclear_and_58_dup_777), .E (
             ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_2__dup_30 (.Q (ENCR_DEV_encry_cnt[2]), .D (
             sclear_and_2_dup_116), .E (ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int
             ), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_1__dup_31 (.Q (ENCR_DEV_encry_cnt[1]), .D (
             sclear_and_1_dup_115), .E (ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int
             ), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_6__dup_26 (.Q (ENCR_DEV_encry_cnt[6]), .D (
             sclear_and_6_dup_120), .E (ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int
             ), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_5__dup_27 (.Q (ENCR_DEV_encry_cnt[5]), .D (
             sclear_and_5_dup_119), .E (ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int
             ), .CLR (RST_int)) ;
    DFN1C0 reg_q_8_ (.Q (ENCR_DEV_cnt_init[8]), .D (sclear_and_8_dup_155), .CLK (
           CLK_int), .CLR (RST_int)) ;
    DFN1C0 reg_q_7_ (.Q (ENCR_DEV_cnt_init[7]), .D (sclear_and_7_dup_154), .CLK (
           CLK_int), .CLR (RST_int)) ;
    DFN1C0 reg_q_9_ (.Q (ENCR_DEV_cnt_init[9]), .D (sclear_and_9_dup_156), .CLK (
           CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_61_ (.Q (ENCR_DEV_reg_str_2[61]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[61]), .E (nx19668z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_58_ (.Q (ENCR_DEV_reg_str_3[58]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[58]), .E (NOT_ENCR_DEV_rtlc15n968__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_62_ (.Q (ENCR_DEV_reg_str_2[62]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[62]), .E (nx19668z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_104_ (.Q (ENCR_DEV_reg_str_3[104]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[104]), .E (
             NOT_ENCR_DEV_rtlc15n968__repl4), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_63_ (.Q (ENCR_DEV_reg_str_2[63]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[63]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_60_ (.Q (ENCR_DEV_reg_str_3[60]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[60]), .E (NOT_ENCR_DEV_rtlc15n968__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_61_ (.Q (ENCR_DEV_reg_str_3[61]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[61]), .E (NOT_ENCR_DEV_rtlc15n968__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_64_ (.Q (ENCR_DEV_reg_str_2[64]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[64]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_62_ (.Q (ENCR_DEV_reg_str_3[62]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[62]), .E (NOT_ENCR_DEV_rtlc15n968__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_65_ (.Q (ENCR_DEV_reg_str_2[65]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[65]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_63_ (.Q (ENCR_DEV_reg_str_3[63]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[63]), .E (NOT_ENCR_DEV_rtlc15n968__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_66_ (.Q (ENCR_DEV_reg_str_2[66]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[66]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_64_ (.Q (ENCR_DEV_reg_str_3[64]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[64]), .E (NOT_ENCR_DEV_rtlc15n968__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_67_ (.Q (ENCR_DEV_reg_str_2[67]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[67]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_92_ (.Q (ENCR_DEV_reg_str_1[92]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[92]), .E (NOT_ENCR_DEV_rtlc15n968__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_110_ (.Q (ENCR_DEV_reg_str_3[110]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[110]), .E (
             NOT_ENCR_DEV_rtlc15n971__repl5), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_25_ (.Q (ENCR_DEV_err_cnt[25]), .D (sclear_and_25_dup_744), .E (
             ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_24_ (.Q (ENCR_DEV_err_cnt[24]), .D (sclear_and_24_dup_743), .E (
             ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_29_ (.Q (ENCR_DEV_err_cnt[29]), .D (sclear_and_29_dup_748), .E (
             ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_28_ (.Q (ENCR_DEV_err_cnt[28]), .D (sclear_and_28_dup_747), .E (
             ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_33_ (.Q (ENCR_DEV_err_cnt[33]), .D (sclear_and_33_dup_752), .E (
             ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_32_ (.Q (ENCR_DEV_err_cnt[32]), .D (sclear_and_32_dup_751), .E (
             ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_37_ (.Q (ENCR_DEV_err_cnt[37]), .D (sclear_and_37_dup_756), .E (
             ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_36_ (.Q (ENCR_DEV_err_cnt[36]), .D (sclear_and_36_dup_755), .E (
             ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_41_ (.Q (ENCR_DEV_err_cnt[41]), .D (sclear_and_41_dup_760), .E (
             ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_40_ (.Q (ENCR_DEV_err_cnt[40]), .D (sclear_and_40_dup_759), .E (
             ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_45_ (.Q (ENCR_DEV_err_cnt[45]), .D (sclear_and_45_dup_764), .E (
             ENCR_DEV_rtlcn483__repl1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_44_ (.Q (ENCR_DEV_err_cnt[44]), .D (sclear_and_44_dup_763), .E (
             ENCR_DEV_rtlcn483__repl0), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_9__dup_2 (.Q (ENCR_DEV_err_cnt[9]), .D (sclear_and_9_dup_728)
             , .E (ENCR_DEV_rtlcn483__repl0), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_8__dup_3 (.Q (ENCR_DEV_err_cnt[8]), .D (sclear_and_8_dup_727)
             , .E (ENCR_DEV_rtlcn483__repl0), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_13_ (.Q (ENCR_DEV_err_cnt[13]), .D (sclear_and_13_dup_732), .E (
             ENCR_DEV_rtlcn483__repl0), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_12_ (.Q (ENCR_DEV_err_cnt[12]), .D (sclear_and_12_dup_731), .E (
             ENCR_DEV_rtlcn483__repl0), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_49_ (.Q (ENCR_DEV_err_cnt[49]), .D (sclear_and_49_dup_768), .E (
             ENCR_DEV_rtlcn483__repl0), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_48_ (.Q (ENCR_DEV_err_cnt[48]), .D (sclear_and_48_dup_767), .E (
             ENCR_DEV_rtlcn483__repl0), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_53_ (.Q (ENCR_DEV_err_cnt[53]), .D (sclear_and_53_dup_772), .E (
             ENCR_DEV_rtlcn483__repl0), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_52_ (.Q (ENCR_DEV_err_cnt[52]), .D (sclear_and_52_dup_771), .E (
             ENCR_DEV_rtlcn483__repl0), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_57_ (.Q (ENCR_DEV_err_cnt[57]), .D (sclear_and_57_dup_776), .E (
             ENCR_DEV_rtlcn483__repl0), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 reg_q_56_ (.Q (ENCR_DEV_err_cnt[56]), .D (sclear_and_56_dup_775), .E (
             ENCR_DEV_rtlcn483__repl0), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 reg_q_4_ (.Q (ENCR_DEV_cnt_init[4]), .D (sclear_and_4_dup_151), .CLK (
           CLK_int), .CLR (RST_int)) ;
    DFN1C0 reg_q_2_ (.Q (ENCR_DEV_cnt_init[2]), .D (sclear_and_2_dup_149), .CLK (
           CLK_int), .CLR (RST_int)) ;
    DFN1C0 reg_q_5_ (.Q (ENCR_DEV_cnt_init[5]), .D (sclear_and_5_dup_152), .CLK (
           CLK_int), .CLR (RST_int)) ;
    DFN1C0 reg_q_1_ (.Q (ENCR_DEV_cnt_init[1]), .D (sclear_and_1_dup_148), .CLK (
           CLK_int), .CLR (RST_int)) ;
    DFN1C0 reg_q_3_ (.Q (ENCR_DEV_cnt_init[3]), .D (sclear_and_3_dup_150), .CLK (
           CLK_int), .CLR (RST_int)) ;
    DFN1C0 reg_q_0_ (.Q (ENCR_DEV_cnt_init[0]), .D (sclear_and_0_dup_147), .CLK (
           CLK_int), .CLR (RST_int)) ;
    DFN1C0 reg_q_6_ (.Q (ENCR_DEV_cnt_init[6]), .D (sclear_and_6_dup_153), .CLK (
           CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_50_ (.Q (ENCR_DEV_reg_str_1[50]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[50]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_57_ (.Q (ENCR_DEV_reg_str_1[57]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[57]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_60_ (.Q (ENCR_DEV_key_reg[60]), .D (
             ENCR_DEV_key_reg_12n5ss1[60]), .E (nx7969z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_95_ (.Q (ENCR_DEV_reg_str_3[95]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[95]), .E (NOT_ENCR_DEV_rtlc15n968__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_102_ (.Q (ENCR_DEV_reg_str_3[102]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[102]), .E (
             NOT_ENCR_DEV_rtlc15n968__repl4), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_77_ (.Q (ENCR_DEV_reg_str_1[77]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[77]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_84_ (.Q (ENCR_DEV_reg_str_1[84]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[84]), .E (NOT_ENCR_DEV_rtlc15n968__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_75_ (.Q (ENCR_DEV_reg_str_2[75]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[75]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_51_ (.Q (ENCR_DEV_reg_str_1[51]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[51]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_61_ (.Q (ENCR_DEV_key_reg[61]), .D (
             ENCR_DEV_key_reg_12n5ss1[61]), .E (nx7969z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_51_ (.Q (ENCR_DEV_reg_str_3[51]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[51]), .E (NOT_ENCR_DEV_rtlc15n968__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_78_ (.Q (ENCR_DEV_reg_str_1[78]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[78]), .E (NOT_ENCR_DEV_rtlc15n968__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_69_ (.Q (ENCR_DEV_reg_str_2[69]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[69]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_52_ (.Q (ENCR_DEV_reg_str_1[52]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[52]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_62_ (.Q (ENCR_DEV_key_reg[62]), .D (
             ENCR_DEV_key_reg_12n5ss1[62]), .E (nx7969z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_97_ (.Q (ENCR_DEV_reg_str_3[97]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[97]), .E (NOT_ENCR_DEV_rtlc15n968__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_79_ (.Q (ENCR_DEV_reg_str_1[79]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[79]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_70_ (.Q (ENCR_DEV_reg_str_2[70]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[70]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_53_ (.Q (ENCR_DEV_reg_str_1[53]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[53]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_63_ (.Q (ENCR_DEV_key_reg[63]), .D (
             ENCR_DEV_key_reg_12n5ss1[63]), .E (nx7969z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_80_ (.Q (ENCR_DEV_reg_str_1[80]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[80]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_71_ (.Q (ENCR_DEV_reg_str_2[71]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[71]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_98_ (.Q (ENCR_DEV_reg_str_3[98]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[98]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_54_ (.Q (ENCR_DEV_reg_str_1[54]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[54]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_64_ (.Q (ENCR_DEV_key_reg[64]), .D (
             ENCR_DEV_key_reg_12n5ss1[64]), .E (nx7969z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_81_ (.Q (ENCR_DEV_reg_str_1[81]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[81]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_72_ (.Q (ENCR_DEV_reg_str_2[72]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[72]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_99_ (.Q (ENCR_DEV_reg_str_3[99]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[99]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_55_ (.Q (ENCR_DEV_reg_str_1[55]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[55]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_65_ (.Q (ENCR_DEV_key_reg[65]), .D (
             ENCR_DEV_key_reg_12n5ss1[65]), .E (nx7969z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_100_ (.Q (ENCR_DEV_reg_str_3[100]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[100]), .E (
             NOT_ENCR_DEV_rtlc15n968__repl3), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_82_ (.Q (ENCR_DEV_reg_str_1[82]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[82]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_73_ (.Q (ENCR_DEV_reg_str_2[73]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[73]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_56_ (.Q (ENCR_DEV_reg_str_1[56]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[56]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_66_ (.Q (ENCR_DEV_key_reg[66]), .D (
             ENCR_DEV_key_reg_12n5ss1[66]), .E (nx7969z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_101_ (.Q (ENCR_DEV_reg_str_3[101]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[101]), .E (
             NOT_ENCR_DEV_rtlc15n968__repl3), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_83_ (.Q (ENCR_DEV_reg_str_1[83]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[83]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_74_ (.Q (ENCR_DEV_reg_str_2[74]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[74]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_60_ (.Q (ENCR_DEV_reg_str_2[60]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[60]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_57_ (.Q (ENCR_DEV_reg_str_3[57]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[57]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_67_ (.Q (ENCR_DEV_key_reg[67]), .D (
             ENCR_DEV_key_reg_12n5ss1[67]), .E (nx7969z1), .CLK (CLK_int), .CLR (
             RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_53_ (.Q (ENCR_DEV_reg_str_2[53]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[53]), .E (NOT_ENCR_DEV_rtlc15n971__repl5
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_50_ (.Q (ENCR_DEV_reg_str_3[50]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[50]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_54_ (.Q (ENCR_DEV_reg_str_2[54]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[54]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_96_ (.Q (ENCR_DEV_reg_str_3[96]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[96]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_55_ (.Q (ENCR_DEV_reg_str_2[55]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[55]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_52_ (.Q (ENCR_DEV_reg_str_3[52]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[52]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_53_ (.Q (ENCR_DEV_reg_str_3[53]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[53]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_56_ (.Q (ENCR_DEV_reg_str_2[56]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[56]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_54_ (.Q (ENCR_DEV_reg_str_3[54]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[54]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_57_ (.Q (ENCR_DEV_reg_str_2[57]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[57]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_55_ (.Q (ENCR_DEV_reg_str_3[55]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[55]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_58_ (.Q (ENCR_DEV_reg_str_2[58]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[58]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_56_ (.Q (ENCR_DEV_reg_str_3[56]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[56]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_59_ (.Q (ENCR_DEV_reg_str_2[59]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[59]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_59_ (.Q (ENCR_DEV_key_reg[59]), .D (
             ENCR_DEV_key_reg_12n5ss1[59]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_42_ (.Q (ENCR_DEV_reg_str_1[42]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[42]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_49_ (.Q (ENCR_DEV_reg_str_1[49]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[49]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_52_ (.Q (ENCR_DEV_key_reg[52]), .D (
             ENCR_DEV_key_reg_12n5ss1[52]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_87_ (.Q (ENCR_DEV_reg_str_3[87]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[87]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_94_ (.Q (ENCR_DEV_reg_str_3[94]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[94]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_69_ (.Q (ENCR_DEV_reg_str_1[69]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[69]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_76_ (.Q (ENCR_DEV_reg_str_1[76]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[76]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_79_ (.Q (ENCR_DEV_key_reg[79]), .D (
             ENCR_DEV_key_reg_12n5ss1[79]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_43_ (.Q (ENCR_DEV_reg_str_1[43]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[43]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_53_ (.Q (ENCR_DEV_key_reg[53]), .D (
             ENCR_DEV_key_reg_12n5ss1[53]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_43_ (.Q (ENCR_DEV_reg_str_3[43]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[43]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_70_ (.Q (ENCR_DEV_reg_str_1[70]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[70]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_44_ (.Q (ENCR_DEV_reg_str_1[44]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[44]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_54_ (.Q (ENCR_DEV_key_reg[54]), .D (
             ENCR_DEV_key_reg_12n5ss1[54]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_89_ (.Q (ENCR_DEV_reg_str_3[89]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[89]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_71_ (.Q (ENCR_DEV_reg_str_1[71]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[71]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_45_ (.Q (ENCR_DEV_reg_str_1[45]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[45]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_55_ (.Q (ENCR_DEV_key_reg[55]), .D (
             ENCR_DEV_key_reg_12n5ss1[55]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_72_ (.Q (ENCR_DEV_reg_str_1[72]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[72]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_90_ (.Q (ENCR_DEV_reg_str_3[90]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[90]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_46_ (.Q (ENCR_DEV_reg_str_1[46]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[46]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_56_ (.Q (ENCR_DEV_key_reg[56]), .D (
             ENCR_DEV_key_reg_12n5ss1[56]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_73_ (.Q (ENCR_DEV_reg_str_1[73]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[73]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_91_ (.Q (ENCR_DEV_reg_str_3[91]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[91]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_47_ (.Q (ENCR_DEV_reg_str_1[47]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[47]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_57_ (.Q (ENCR_DEV_key_reg[57]), .D (
             ENCR_DEV_key_reg_12n5ss1[57]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_92_ (.Q (ENCR_DEV_reg_str_3[92]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[92]), .E (NOT_ENCR_DEV_rtlc15n968__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_74_ (.Q (ENCR_DEV_reg_str_1[74]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[74]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_48_ (.Q (ENCR_DEV_reg_str_1[48]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[48]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_58_ (.Q (ENCR_DEV_key_reg[58]), .D (
             ENCR_DEV_key_reg_12n5ss1[58]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_93_ (.Q (ENCR_DEV_reg_str_3[93]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[93]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_75_ (.Q (ENCR_DEV_reg_str_1[75]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[75]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_52_ (.Q (ENCR_DEV_reg_str_2[52]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[52]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_49_ (.Q (ENCR_DEV_reg_str_3[49]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[49]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_45_ (.Q (ENCR_DEV_reg_str_2[45]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[45]), .E (NOT_ENCR_DEV_rtlc15n971__repl4
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_42_ (.Q (ENCR_DEV_reg_str_3[42]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[42]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_46_ (.Q (ENCR_DEV_reg_str_2[46]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[46]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_88_ (.Q (ENCR_DEV_reg_str_3[88]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[88]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_47_ (.Q (ENCR_DEV_reg_str_2[47]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[47]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_44_ (.Q (ENCR_DEV_reg_str_3[44]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[44]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_45_ (.Q (ENCR_DEV_reg_str_3[45]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[45]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_48_ (.Q (ENCR_DEV_reg_str_2[48]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[48]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_46_ (.Q (ENCR_DEV_reg_str_3[46]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[46]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_49_ (.Q (ENCR_DEV_reg_str_2[49]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[49]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_47_ (.Q (ENCR_DEV_reg_str_3[47]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[47]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_50_ (.Q (ENCR_DEV_reg_str_2[50]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[50]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_48_ (.Q (ENCR_DEV_reg_str_3[48]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[48]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_51_ (.Q (ENCR_DEV_reg_str_2[51]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[51]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_51_ (.Q (ENCR_DEV_key_reg[51]), .D (
             ENCR_DEV_key_reg_12n5ss1[51]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_78_ (.Q (ENCR_DEV_key_reg[78]), .D (
             ENCR_DEV_key_reg_12n5ss1[78]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_34_ (.Q (ENCR_DEV_reg_str_1[34]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[34]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_41_ (.Q (ENCR_DEV_reg_str_1[41]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[41]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_44_ (.Q (ENCR_DEV_key_reg[44]), .D (
             ENCR_DEV_key_reg_12n5ss1[44]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_79_ (.Q (ENCR_DEV_reg_str_3[79]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[79]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_86_ (.Q (ENCR_DEV_reg_str_3[86]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[86]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_68_ (.Q (ENCR_DEV_reg_str_1[68]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[68]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_71_ (.Q (ENCR_DEV_key_reg[71]), .D (
             ENCR_DEV_key_reg_12n5ss1[71]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_35_ (.Q (ENCR_DEV_reg_str_1[35]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[35]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_45_ (.Q (ENCR_DEV_key_reg[45]), .D (
             ENCR_DEV_key_reg_12n5ss1[45]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_35_ (.Q (ENCR_DEV_reg_str_3[35]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[35]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_72_ (.Q (ENCR_DEV_key_reg[72]), .D (
             ENCR_DEV_key_reg_12n5ss1[72]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_36_ (.Q (ENCR_DEV_reg_str_1[36]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[36]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_46_ (.Q (ENCR_DEV_key_reg[46]), .D (
             ENCR_DEV_key_reg_12n5ss1[46]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_81_ (.Q (ENCR_DEV_reg_str_3[81]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[81]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_73_ (.Q (ENCR_DEV_key_reg[73]), .D (
             ENCR_DEV_key_reg_12n5ss1[73]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_37_ (.Q (ENCR_DEV_reg_str_1[37]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[37]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_47_ (.Q (ENCR_DEV_key_reg[47]), .D (
             ENCR_DEV_key_reg_12n5ss1[47]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_74_ (.Q (ENCR_DEV_key_reg[74]), .D (
             ENCR_DEV_key_reg_12n5ss1[74]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_82_ (.Q (ENCR_DEV_reg_str_3[82]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[82]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_38_ (.Q (ENCR_DEV_reg_str_1[38]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[38]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_48_ (.Q (ENCR_DEV_key_reg[48]), .D (
             ENCR_DEV_key_reg_12n5ss1[48]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_75_ (.Q (ENCR_DEV_key_reg[75]), .D (
             ENCR_DEV_key_reg_12n5ss1[75]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_83_ (.Q (ENCR_DEV_reg_str_3[83]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[83]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_39_ (.Q (ENCR_DEV_reg_str_1[39]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[39]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_49_ (.Q (ENCR_DEV_key_reg[49]), .D (
             ENCR_DEV_key_reg_12n5ss1[49]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_84_ (.Q (ENCR_DEV_reg_str_3[84]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[84]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_66_ (.Q (ENCR_DEV_reg_str_1[66]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[66]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_76_ (.Q (ENCR_DEV_key_reg[76]), .D (
             ENCR_DEV_key_reg_12n5ss1[76]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_40_ (.Q (ENCR_DEV_reg_str_1[40]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[40]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_50_ (.Q (ENCR_DEV_key_reg[50]), .D (
             ENCR_DEV_key_reg_12n5ss1[50]), .E (NOT_ENCR_DEV_rtlc12n435__repl2)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_85_ (.Q (ENCR_DEV_reg_str_3[85]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[85]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_67_ (.Q (ENCR_DEV_reg_str_1[67]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[67]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_77_ (.Q (ENCR_DEV_key_reg[77]), .D (
             ENCR_DEV_key_reg_12n5ss1[77]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_44_ (.Q (ENCR_DEV_reg_str_2[44]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[44]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_41_ (.Q (ENCR_DEV_reg_str_3[41]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[41]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_37_ (.Q (ENCR_DEV_reg_str_2[37]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[37]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_34_ (.Q (ENCR_DEV_reg_str_3[34]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[34]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_38_ (.Q (ENCR_DEV_reg_str_2[38]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[38]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_80_ (.Q (ENCR_DEV_reg_str_3[80]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[80]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_39_ (.Q (ENCR_DEV_reg_str_2[39]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[39]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_36_ (.Q (ENCR_DEV_reg_str_3[36]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[36]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_37_ (.Q (ENCR_DEV_reg_str_3[37]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[37]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_40_ (.Q (ENCR_DEV_reg_str_2[40]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[40]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_38_ (.Q (ENCR_DEV_reg_str_3[38]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[38]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_41_ (.Q (ENCR_DEV_reg_str_2[41]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[41]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_39_ (.Q (ENCR_DEV_reg_str_3[39]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[39]), .E (NOT_ENCR_DEV_rtlc15n968__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_42_ (.Q (ENCR_DEV_reg_str_2[42]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[42]), .E (NOT_ENCR_DEV_rtlc15n971__repl3
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_40_ (.Q (ENCR_DEV_reg_str_3[40]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[40]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_43_ (.Q (ENCR_DEV_reg_str_2[43]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[43]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_43_ (.Q (ENCR_DEV_key_reg[43]), .D (
             ENCR_DEV_key_reg_12n5ss1[43]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_70_ (.Q (ENCR_DEV_key_reg[70]), .D (
             ENCR_DEV_key_reg_12n5ss1[70]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_26_ (.Q (ENCR_DEV_reg_str_1[26]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[26]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_33_ (.Q (ENCR_DEV_reg_str_1[33]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[33]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_36_ (.Q (ENCR_DEV_key_reg[36]), .D (
             ENCR_DEV_key_reg_12n5ss1[36]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_71_ (.Q (ENCR_DEV_reg_str_3[71]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[71]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_78_ (.Q (ENCR_DEV_reg_str_3[78]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[78]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_27_ (.Q (ENCR_DEV_reg_str_1[27]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[27]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_37_ (.Q (ENCR_DEV_key_reg[37]), .D (
             ENCR_DEV_key_reg_12n5ss1[37]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_27_ (.Q (ENCR_DEV_reg_str_3[27]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[27]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_28_ (.Q (ENCR_DEV_reg_str_1[28]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[28]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_38_ (.Q (ENCR_DEV_key_reg[38]), .D (
             ENCR_DEV_key_reg_12n5ss1[38]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_73_ (.Q (ENCR_DEV_reg_str_3[73]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[73]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_29_ (.Q (ENCR_DEV_reg_str_1[29]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[29]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_39_ (.Q (ENCR_DEV_key_reg[39]), .D (
             ENCR_DEV_key_reg_12n5ss1[39]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_74_ (.Q (ENCR_DEV_reg_str_3[74]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[74]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_30_ (.Q (ENCR_DEV_reg_str_1[30]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[30]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_40_ (.Q (ENCR_DEV_key_reg[40]), .D (
             ENCR_DEV_key_reg_12n5ss1[40]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_75_ (.Q (ENCR_DEV_reg_str_3[75]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[75]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_31_ (.Q (ENCR_DEV_reg_str_1[31]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[31]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_41_ (.Q (ENCR_DEV_key_reg[41]), .D (
             ENCR_DEV_key_reg_12n5ss1[41]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_76_ (.Q (ENCR_DEV_reg_str_3[76]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[76]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_68_ (.Q (ENCR_DEV_key_reg[68]), .D (
             ENCR_DEV_key_reg_12n5ss1[68]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_32_ (.Q (ENCR_DEV_reg_str_1[32]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[32]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_42_ (.Q (ENCR_DEV_key_reg[42]), .D (
             ENCR_DEV_key_reg_12n5ss1[42]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_77_ (.Q (ENCR_DEV_reg_str_3[77]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[77]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_69_ (.Q (ENCR_DEV_key_reg[69]), .D (
             ENCR_DEV_key_reg_12n5ss1[69]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_36_ (.Q (ENCR_DEV_reg_str_2[36]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[36]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_33_ (.Q (ENCR_DEV_reg_str_3[33]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[33]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_29_ (.Q (ENCR_DEV_reg_str_2[29]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[29]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_26_ (.Q (ENCR_DEV_reg_str_3[26]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[26]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_30_ (.Q (ENCR_DEV_reg_str_2[30]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[30]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_72_ (.Q (ENCR_DEV_reg_str_3[72]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[72]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_31_ (.Q (ENCR_DEV_reg_str_2[31]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[31]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_28_ (.Q (ENCR_DEV_reg_str_3[28]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[28]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_29_ (.Q (ENCR_DEV_reg_str_3[29]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[29]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_32_ (.Q (ENCR_DEV_reg_str_2[32]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[32]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_30_ (.Q (ENCR_DEV_reg_str_3[30]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[30]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_33_ (.Q (ENCR_DEV_reg_str_2[33]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[33]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_31_ (.Q (ENCR_DEV_reg_str_3[31]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[31]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_34_ (.Q (ENCR_DEV_reg_str_2[34]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[34]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_32_ (.Q (ENCR_DEV_reg_str_3[32]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[32]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_35_ (.Q (ENCR_DEV_reg_str_2[35]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[35]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_35_ (.Q (ENCR_DEV_key_reg[35]), .D (
             ENCR_DEV_key_reg_12n5ss1[35]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_18_ (.Q (ENCR_DEV_reg_str_1[18]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[18]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_25_ (.Q (ENCR_DEV_reg_str_1[25]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[25]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_28_ (.Q (ENCR_DEV_key_reg[28]), .D (
             ENCR_DEV_key_reg_12n5ss1[28]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_70_ (.Q (ENCR_DEV_reg_str_3[70]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[70]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_19_ (.Q (ENCR_DEV_reg_str_1[19]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[19]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_29_ (.Q (ENCR_DEV_key_reg[29]), .D (
             ENCR_DEV_key_reg_12n5ss1[29]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_19_ (.Q (ENCR_DEV_reg_str_3[19]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[19]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_20_ (.Q (ENCR_DEV_reg_str_1[20]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[20]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_30_ (.Q (ENCR_DEV_key_reg[30]), .D (
             ENCR_DEV_key_reg_12n5ss1[30]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_21_ (.Q (ENCR_DEV_reg_str_1[21]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[21]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_31_ (.Q (ENCR_DEV_key_reg[31]), .D (
             ENCR_DEV_key_reg_12n5ss1[31]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_66_ (.Q (ENCR_DEV_reg_str_3[66]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[66]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_22_ (.Q (ENCR_DEV_reg_str_1[22]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[22]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_32_ (.Q (ENCR_DEV_key_reg[32]), .D (
             ENCR_DEV_key_reg_12n5ss1[32]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_67_ (.Q (ENCR_DEV_reg_str_3[67]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[67]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_23_ (.Q (ENCR_DEV_reg_str_1[23]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[23]), .E (NOT_ENCR_DEV_rtlc15n971__repl2
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_33_ (.Q (ENCR_DEV_key_reg[33]), .D (
             ENCR_DEV_key_reg_12n5ss1[33]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_68_ (.Q (ENCR_DEV_reg_str_3[68]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[68]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_24_ (.Q (ENCR_DEV_reg_str_1[24]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[24]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_34_ (.Q (ENCR_DEV_key_reg[34]), .D (
             ENCR_DEV_key_reg_12n5ss1[34]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_69_ (.Q (ENCR_DEV_reg_str_3[69]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[69]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_28_ (.Q (ENCR_DEV_reg_str_2[28]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[28]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_25_ (.Q (ENCR_DEV_reg_str_3[25]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[25]), .E (NOT_ENCR_DEV_rtlc15n968__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_21_ (.Q (ENCR_DEV_reg_str_2[21]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[21]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_18_ (.Q (ENCR_DEV_reg_str_3[18]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[18]), .E (NOT_ENCR_DEV_rtlc15n968__repl0
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_22_ (.Q (ENCR_DEV_reg_str_2[22]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[22]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_23_ (.Q (ENCR_DEV_reg_str_2[23]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[23]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_20_ (.Q (ENCR_DEV_reg_str_3[20]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[20]), .E (NOT_ENCR_DEV_rtlc15n968__repl0
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_21_ (.Q (ENCR_DEV_reg_str_3[21]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[21]), .E (NOT_ENCR_DEV_rtlc15n968__repl0
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_24_ (.Q (ENCR_DEV_reg_str_2[24]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[24]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_22_ (.Q (ENCR_DEV_reg_str_3[22]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[22]), .E (NOT_ENCR_DEV_rtlc15n968__repl0
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_25_ (.Q (ENCR_DEV_reg_str_2[25]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[25]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_23_ (.Q (ENCR_DEV_reg_str_3[23]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[23]), .E (NOT_ENCR_DEV_rtlc15n968__repl0
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_26_ (.Q (ENCR_DEV_reg_str_2[26]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[26]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_24_ (.Q (ENCR_DEV_reg_str_3[24]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[24]), .E (NOT_ENCR_DEV_rtlc15n968__repl0
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_27_ (.Q (ENCR_DEV_reg_str_2[27]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[27]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_27_ (.Q (ENCR_DEV_key_reg[27]), .D (
             ENCR_DEV_key_reg_12n5ss1[27]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_10_ (.Q (ENCR_DEV_reg_str_1[10]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[10]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_17_ (.Q (ENCR_DEV_reg_str_1[17]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[17]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_20_ (.Q (ENCR_DEV_key_reg[20]), .D (
             ENCR_DEV_key_reg_12n5ss1[20]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_11_ (.Q (ENCR_DEV_reg_str_1[11]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[11]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_21_ (.Q (ENCR_DEV_key_reg[21]), .D (
             ENCR_DEV_key_reg_12n5ss1[21]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_11_ (.Q (ENCR_DEV_reg_str_3[11]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[11]), .E (NOT_ENCR_DEV_rtlc15n968__repl0
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_12_ (.Q (ENCR_DEV_reg_str_1[12]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[12]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_22_ (.Q (ENCR_DEV_key_reg[22]), .D (
             ENCR_DEV_key_reg_12n5ss1[22]), .E (NOT_ENCR_DEV_rtlc12n435__repl1)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_13_ (.Q (ENCR_DEV_reg_str_1[13]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[13]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_23_ (.Q (ENCR_DEV_key_reg[23]), .D (
             ENCR_DEV_key_reg_12n5ss1[23]), .E (NOT_ENCR_DEV_rtlc12n435__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_14_ (.Q (ENCR_DEV_reg_str_1[14]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[14]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_24_ (.Q (ENCR_DEV_key_reg[24]), .D (
             ENCR_DEV_key_reg_12n5ss1[24]), .E (NOT_ENCR_DEV_rtlc12n435__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_15_ (.Q (ENCR_DEV_reg_str_1[15]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[15]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_25_ (.Q (ENCR_DEV_key_reg[25]), .D (
             ENCR_DEV_key_reg_12n5ss1[25]), .E (NOT_ENCR_DEV_rtlc12n435__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_16_ (.Q (ENCR_DEV_reg_str_1[16]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[16]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_26_ (.Q (ENCR_DEV_key_reg[26]), .D (
             ENCR_DEV_key_reg_12n5ss1[26]), .E (NOT_ENCR_DEV_rtlc12n435__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_20_ (.Q (ENCR_DEV_reg_str_2[20]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[20]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_17_ (.Q (ENCR_DEV_reg_str_3[17]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[17]), .E (NOT_ENCR_DEV_rtlc15n968__repl0
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_13_ (.Q (ENCR_DEV_reg_str_2[13]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[13]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_10_ (.Q (ENCR_DEV_reg_str_3[10]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[10]), .E (NOT_ENCR_DEV_rtlc15n968__repl0
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_14_ (.Q (ENCR_DEV_reg_str_2[14]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[14]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_15_ (.Q (ENCR_DEV_reg_str_2[15]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[15]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_12_ (.Q (ENCR_DEV_reg_str_3[12]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[12]), .E (NOT_ENCR_DEV_rtlc15n968__repl0
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_13_ (.Q (ENCR_DEV_reg_str_3[13]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[13]), .E (NOT_ENCR_DEV_rtlc15n968__repl0
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_16_ (.Q (ENCR_DEV_reg_str_2[16]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[16]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_14_ (.Q (ENCR_DEV_reg_str_3[14]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[14]), .E (NOT_ENCR_DEV_rtlc15n968__repl0
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_17_ (.Q (ENCR_DEV_reg_str_2[17]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[17]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_15_ (.Q (ENCR_DEV_reg_str_3[15]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[15]), .E (NOT_ENCR_DEV_rtlc15n968__repl0
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_18_ (.Q (ENCR_DEV_reg_str_2[18]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[18]), .E (NOT_ENCR_DEV_rtlc15n971__repl1
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_16_ (.Q (ENCR_DEV_reg_str_3[16]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[16]), .E (NOT_ENCR_DEV_rtlc15n968__repl0
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_19_ (.Q (ENCR_DEV_reg_str_2[19]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[19]), .E (NOT_ENCR_DEV_rtlc15n971__repl0
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_19_ (.Q (ENCR_DEV_key_reg[19]), .D (
             ENCR_DEV_key_reg_12n5ss1[19]), .E (NOT_ENCR_DEV_rtlc12n435__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_2_ (.Q (ENCR_DEV_reg_str_1[2]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[2]), .E (NOT_ENCR_DEV_rtlc15n971__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_9_ (.Q (ENCR_DEV_reg_str_1[9]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[9]), .E (NOT_ENCR_DEV_rtlc15n971__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_12_ (.Q (ENCR_DEV_key_reg[12]), .D (
             ENCR_DEV_key_reg_12n5ss1[12]), .E (NOT_ENCR_DEV_rtlc12n435__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_3_ (.Q (ENCR_DEV_reg_str_1[3]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[3]), .E (NOT_ENCR_DEV_rtlc15n971__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_13_ (.Q (ENCR_DEV_key_reg[13]), .D (
             ENCR_DEV_key_reg_12n5ss1[13]), .E (NOT_ENCR_DEV_rtlc12n435__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_3_ (.Q (ENCR_DEV_reg_str_3[3]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[3]), .E (NOT_ENCR_DEV_rtlc15n968__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_4_ (.Q (ENCR_DEV_reg_str_1[4]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[4]), .E (NOT_ENCR_DEV_rtlc15n971__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_14_ (.Q (ENCR_DEV_key_reg[14]), .D (
             ENCR_DEV_key_reg_12n5ss1[14]), .E (NOT_ENCR_DEV_rtlc12n435__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_5_ (.Q (ENCR_DEV_reg_str_1[5]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[5]), .E (NOT_ENCR_DEV_rtlc15n971__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_15_ (.Q (ENCR_DEV_key_reg[15]), .D (
             ENCR_DEV_key_reg_12n5ss1[15]), .E (NOT_ENCR_DEV_rtlc12n435__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_6_ (.Q (ENCR_DEV_reg_str_1[6]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[6]), .E (NOT_ENCR_DEV_rtlc15n971__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_16_ (.Q (ENCR_DEV_key_reg[16]), .D (
             ENCR_DEV_key_reg_12n5ss1[16]), .E (NOT_ENCR_DEV_rtlc12n435__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_7_ (.Q (ENCR_DEV_reg_str_1[7]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[7]), .E (NOT_ENCR_DEV_rtlc15n971__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_17_ (.Q (ENCR_DEV_key_reg[17]), .D (
             ENCR_DEV_key_reg_12n5ss1[17]), .E (NOT_ENCR_DEV_rtlc12n435__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_8_ (.Q (ENCR_DEV_reg_str_1[8]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[8]), .E (NOT_ENCR_DEV_rtlc15n971__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_18_ (.Q (ENCR_DEV_key_reg[18]), .D (
             ENCR_DEV_key_reg_12n5ss1[18]), .E (NOT_ENCR_DEV_rtlc12n435__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_12_ (.Q (ENCR_DEV_reg_str_2[12]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[12]), .E (NOT_ENCR_DEV_rtlc15n971__repl0
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_9_ (.Q (ENCR_DEV_reg_str_3[9]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[9]), .E (NOT_ENCR_DEV_rtlc15n968__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_5_ (.Q (ENCR_DEV_reg_str_2[5]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[5]), .E (NOT_ENCR_DEV_rtlc15n971__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_2_ (.Q (ENCR_DEV_reg_str_3[2]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[2]), .E (NOT_ENCR_DEV_rtlc15n968__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_6_ (.Q (ENCR_DEV_reg_str_2[6]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[6]), .E (NOT_ENCR_DEV_rtlc15n971__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_7_ (.Q (ENCR_DEV_reg_str_2[7]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[7]), .E (NOT_ENCR_DEV_rtlc15n971__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_4_ (.Q (ENCR_DEV_reg_str_3[4]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[4]), .E (NOT_ENCR_DEV_rtlc15n968__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_5_ (.Q (ENCR_DEV_reg_str_3[5]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[5]), .E (NOT_ENCR_DEV_rtlc15n968__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_8_ (.Q (ENCR_DEV_reg_str_2[8]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[8]), .E (NOT_ENCR_DEV_rtlc15n971__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_6_ (.Q (ENCR_DEV_reg_str_3[6]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[6]), .E (NOT_ENCR_DEV_rtlc15n968__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_9_ (.Q (ENCR_DEV_reg_str_2[9]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[9]), .E (NOT_ENCR_DEV_rtlc15n971__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_7_ (.Q (ENCR_DEV_reg_str_3[7]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[7]), .E (NOT_ENCR_DEV_rtlc15n968__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_10_ (.Q (ENCR_DEV_reg_str_2[10]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[10]), .E (NOT_ENCR_DEV_rtlc15n971__repl0
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_8_ (.Q (ENCR_DEV_reg_str_3[8]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[8]), .E (NOT_ENCR_DEV_rtlc15n968__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_11_ (.Q (ENCR_DEV_reg_str_2[11]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[11]), .E (NOT_ENCR_DEV_rtlc15n971__repl0
             ), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_11_ (.Q (ENCR_DEV_key_reg[11]), .D (
             ENCR_DEV_key_reg_12n5ss1[11]), .E (NOT_ENCR_DEV_rtlc12n435__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_1_ (.Q (ENCR_DEV_reg_str_1[1]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[1]), .E (NOT_ENCR_DEV_rtlc15n971__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_4_ (.Q (ENCR_DEV_key_reg[4]), .D (
             ENCR_DEV_key_reg_12n5ss1[4]), .E (NOT_ENCR_DEV_rtlc12n435__repl0), 
             .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_5_ (.Q (ENCR_DEV_key_reg[5]), .D (
             ENCR_DEV_key_reg_12n5ss1[5]), .E (NOT_ENCR_DEV_rtlc12n435__repl0), 
             .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_6_ (.Q (ENCR_DEV_key_reg[6]), .D (
             ENCR_DEV_key_reg_12n5ss1[6]), .E (NOT_ENCR_DEV_rtlc12n435__repl0), 
             .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_7_ (.Q (ENCR_DEV_key_reg[7]), .D (
             ENCR_DEV_key_reg_12n5ss1[7]), .E (NOT_ENCR_DEV_rtlc12n435__repl0), 
             .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_8_ (.Q (ENCR_DEV_key_reg[8]), .D (
             ENCR_DEV_key_reg_12n5ss1[8]), .E (NOT_ENCR_DEV_rtlc12n435__repl0), 
             .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_9_ (.Q (ENCR_DEV_key_reg[9]), .D (
             ENCR_DEV_key_reg_12n5ss1[9]), .E (NOT_ENCR_DEV_rtlc12n435__repl0), 
             .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_1_0_ (.Q (ENCR_DEV_reg_str_1[0]), .D (
             ENCR_DEV_reg_str_1_15n2ss1[0]), .E (NOT_ENCR_DEV_rtlc15n971__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_10_ (.Q (ENCR_DEV_key_reg[10]), .D (
             ENCR_DEV_key_reg_12n5ss1[10]), .E (NOT_ENCR_DEV_rtlc12n435__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_4_ (.Q (ENCR_DEV_reg_str_2[4]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[4]), .E (NOT_ENCR_DEV_rtlc15n971__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_1_ (.Q (ENCR_DEV_reg_str_3[1]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[1]), .E (NOT_ENCR_DEV_rtlc15n968__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_0_ (.Q (ENCR_DEV_reg_str_2[0]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[0]), .E (NOT_ENCR_DEV_rtlc15n971__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_1_ (.Q (ENCR_DEV_reg_str_2[1]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[1]), .E (NOT_ENCR_DEV_rtlc15n971__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_2_ (.Q (ENCR_DEV_reg_str_2[2]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[2]), .E (NOT_ENCR_DEV_rtlc15n971__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_3_0_ (.Q (ENCR_DEV_reg_str_3[0]), .D (
             ENCR_DEV_reg_str_3_15n2ss1[0]), .E (NOT_ENCR_DEV_rtlc15n968__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_reg_str_2_3_ (.Q (ENCR_DEV_reg_str_2[3]), .D (
             ENCR_DEV_reg_str_2_15n2ss1[3]), .E (NOT_ENCR_DEV_rtlc15n971__repl0)
             , .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_3_ (.Q (ENCR_DEV_key_reg[3]), .D (
             ENCR_DEV_key_reg_12n5ss1[3]), .E (NOT_ENCR_DEV_rtlc12n435__repl0), 
             .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_2_ (.Q (ENCR_DEV_key_reg[2]), .D (
             ENCR_DEV_key_reg_12n5ss1[2]), .E (NOT_ENCR_DEV_rtlc12n435__repl0), 
             .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_1_ (.Q (ENCR_DEV_key_reg[1]), .D (
             ENCR_DEV_key_reg_12n5ss1[1]), .E (NOT_ENCR_DEV_rtlc12n435__repl0), 
             .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 ENCR_DEV_reg_key_reg_0_ (.Q (ENCR_DEV_key_reg[0]), .D (
             ENCR_DEV_key_reg_12n5ss1[0]), .E (NOT_ENCR_DEV_rtlc12n435__repl0), 
             .CLK (CLK_int), .CLR (RST_int)) ;
    CLKBUF CLK_ibuf (.Y (CLK_int), .PAD (CLK)) ;
    CLKBUF RST_ibuf (.Y (RST_int), .PAD (RST)) ;
    CLKINT buf_ENCR_DEV_prev_6_ (.Y (ENCR_DEV_prev_6__int), .A (ENCR_DEV_prev[6]
           )) ;
    CLKINT buf_NOT_FIFO_DEV_ix32158z56071 (.Y (NOT_FIFO_DEV_rtlc5n43_int), .A (
           nx32158z2)) ;
    CLKINT buf_b_0_ (.Y (b_0__int), .A (b_0_)) ;
    CLKINT buf_NOT_ENCR_DEV_ix37688z56070 (.Y (NOT_ENCR_DEV_rtlcn261_int), .A (
           nx37688z1)) ;
    AO1A NOT_ENCR_DEV_rtlc12n435__repl0_rename1015 (.Y (
         NOT_ENCR_DEV_rtlc12n435__repl0), .A (STB_KEY_int), .B (nx18636z1), .C (
         nx18636z2)) ;
    AO1A NOT_ENCR_DEV_rtlc12n435__repl1_rename1016 (.Y (
         NOT_ENCR_DEV_rtlc12n435__repl1), .A (STB_KEY_int), .B (nx18636z1), .C (
         nx18636z2)) ;
    AO1A NOT_ENCR_DEV_rtlc12n435__repl2_rename1017 (.Y (
         NOT_ENCR_DEV_rtlc12n435__repl2), .A (STB_KEY_int), .B (nx18636z1), .C (
         nx18636z2)) ;
    DFN1E0C0 FIFO_DEV_modgen_counter_rtlc_radd_N1_reg_q_5__dup__repl0 (.Q (
             FIFO_DEV_rtlc_radd_N1_5___repl0), .D (
             FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_5_), .E (nx12521z2), .CLK (
             CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 FIFO_DEV_modgen_counter_rtlc_radd_N1_reg_q_5__dup__repl1 (.Q (
             FIFO_DEV_rtlc_radd_N1_5___repl1), .D (
             FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_5_), .E (nx12521z2), .CLK (
             CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 FIFO_DEV_modgen_counter_rtlc_radd_N1_reg_q_3__dup__repl0 (.Q (
             FIFO_DEV_rtlc_radd_N1_3___repl0), .D (
             FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_3_), .E (nx12521z2), .CLK (
             CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 FIFO_DEV_modgen_counter_rtlc_radd_N1_reg_q_2__dup__repl0 (.Q (
             FIFO_DEV_rtlc_radd_N1_2___repl0), .D (
             FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_2_), .E (nx12521z2), .CLK (
             CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 FIFO_DEV_modgen_counter_rtlc_radd_N1_reg_q_2__dup__repl1 (.Q (
             FIFO_DEV_rtlc_radd_N1_2___repl1), .D (
             FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_2_), .E (nx12521z2), .CLK (
             CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 FIFO_DEV_modgen_counter_rtlc_radd_N1_reg_q_2__dup__repl2 (.Q (
             FIFO_DEV_rtlc_radd_N1_2___repl2), .D (
             FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_2_), .E (nx12521z2), .CLK (
             CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 FIFO_DEV_modgen_counter_rtlc_radd_N1_reg_q_1__dup__repl0 (.Q (
             FIFO_DEV_rtlc_radd_N1_1___repl0), .D (
             FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_1_), .E (nx12521z2), .CLK (
             CLK_int), .CLR (RST_int)) ;
    DFN1E0C0 FIFO_DEV_modgen_counter_rtlc_radd_N1_reg_q_0__dup__repl0 (.Q (
             FIFO_DEV_rtlc_radd_N1_0___repl0), .D (
             FIFO_DEV_modgen_counter_rtlc_radd_N1_inc_d_0_), .E (nx12521z2), .CLK (
             CLK_int), .CLR (RST_int)) ;
    NAND3C NOT_ENCR_DEV_rtlc15n971__repl0_rename1018 (.Y (
           NOT_ENCR_DEV_rtlc15n971__repl0), .A (ENCR_DEV_rtlc15_PS14_n166), .B (
           ENCR_DEV_prev[3]), .C (ENCR_DEV_rtlcn483__repl0)) ;
    NAND3C NOT_ENCR_DEV_rtlc15n971__repl1_rename1019 (.Y (
           NOT_ENCR_DEV_rtlc15n971__repl1), .A (ENCR_DEV_rtlc15_PS14_n166), .B (
           ENCR_DEV_prev[3]), .C (ENCR_DEV_rtlcn483__repl0)) ;
    NAND3C NOT_ENCR_DEV_rtlc15n971__repl2_rename1020 (.Y (
           NOT_ENCR_DEV_rtlc15n971__repl2), .A (ENCR_DEV_rtlc15_PS14_n166), .B (
           ENCR_DEV_prev[3]), .C (ENCR_DEV_rtlcn483__repl0)) ;
    NAND3C NOT_ENCR_DEV_rtlc15n971__repl3_rename1021 (.Y (
           NOT_ENCR_DEV_rtlc15n971__repl3), .A (ENCR_DEV_rtlc15_PS14_n166), .B (
           ENCR_DEV_prev[3]), .C (ENCR_DEV_rtlcn483__repl0)) ;
    NAND3C NOT_ENCR_DEV_rtlc15n971__repl4_rename1022 (.Y (
           NOT_ENCR_DEV_rtlc15n971__repl4), .A (ENCR_DEV_rtlc15_PS14_n166), .B (
           ENCR_DEV_prev[3]), .C (ENCR_DEV_rtlcn483__repl0)) ;
    NAND3C NOT_ENCR_DEV_rtlc15n971__repl5_rename1023 (.Y (
           NOT_ENCR_DEV_rtlc15n971__repl5), .A (ENCR_DEV_rtlc15_PS14_n166), .B (
           ENCR_DEV_prev[3]), .C (ENCR_DEV_rtlcn483__repl0)) ;
    DFN1C0 ENCR_DEV_reg_prev_5___repl0 (.Q (ENCR_DEV_prev_5___repl0), .D (
           nx36622z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_prev_5___repl1 (.Q (ENCR_DEV_prev_5___repl1), .D (
           nx36622z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_prev_5___repl2 (.Q (ENCR_DEV_prev_5___repl2), .D (
           nx36622z1), .CLK (CLK_int), .CLR (RST_int)) ;
    AO1D NOT_ENCR_DEV_rtlc15n968__repl0_rename1024 (.Y (
         NOT_ENCR_DEV_rtlc15n968__repl0), .A (nx23410z1), .B (nx3438z4), .C (
         ENCR_DEV_rtlcn483__repl0)) ;
    AO1D NOT_ENCR_DEV_rtlc15n968__repl1_rename1025 (.Y (
         NOT_ENCR_DEV_rtlc15n968__repl1), .A (nx23410z1), .B (nx3438z4), .C (
         ENCR_DEV_rtlcn483__repl0)) ;
    AO1D NOT_ENCR_DEV_rtlc15n968__repl2_rename1026 (.Y (
         NOT_ENCR_DEV_rtlc15n968__repl2), .A (nx23410z1), .B (nx3438z4), .C (
         ENCR_DEV_rtlcn483__repl0)) ;
    AO1D NOT_ENCR_DEV_rtlc15n968__repl3_rename1027 (.Y (
         NOT_ENCR_DEV_rtlc15n968__repl3), .A (nx23410z1), .B (nx3438z4), .C (
         ENCR_DEV_rtlcn483__repl0)) ;
    AO1D NOT_ENCR_DEV_rtlc15n968__repl4_rename1028 (.Y (
         NOT_ENCR_DEV_rtlc15n968__repl4), .A (nx23410z1), .B (nx3438z4), .C (
         ENCR_DEV_rtlcn483__repl0)) ;
    DFN1C0 ENCR_DEV_reg_prev_1___repl0 (.Q (ENCR_DEV_prev_1___repl0), .D (
           nx3438z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_prev_1___repl1 (.Q (ENCR_DEV_prev_1___repl1), .D (
           nx3438z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_prev_1___repl2 (.Q (ENCR_DEV_prev_1___repl2), .D (
           nx3438z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_prev_1___repl3 (.Q (ENCR_DEV_prev_1___repl3), .D (
           nx3438z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_prev_1___repl4 (.Q (ENCR_DEV_prev_1___repl4), .D (
           nx3438z1), .CLK (CLK_int), .CLR (RST_int)) ;
    AND2A ENCR_DEV_rtlcn483__repl0_rename1029 (.Y (ENCR_DEV_rtlcn483__repl0), .A (
          ENCR_DEV_strob_data_tmp), .B (ENCR_DEV_prev[2])) ;
    AND2A ENCR_DEV_rtlcn483__repl1_rename1030 (.Y (ENCR_DEV_rtlcn483__repl1), .A (
          ENCR_DEV_strob_data_tmp), .B (ENCR_DEV_prev[2])) ;
    AND2A ENCR_DEV_rtlcn483__repl2_rename1031 (.Y (ENCR_DEV_rtlcn483__repl2), .A (
          ENCR_DEV_strob_data_tmp), .B (ENCR_DEV_prev[2])) ;
    DFN1C0 ENCR_DEV_reg_prev_8___repl0 (.Q (ENCR_DEV_prev_8___repl0), .D (
           nx15492z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_prev_8___repl1 (.Q (ENCR_DEV_prev_8___repl1), .D (
           nx15492z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_prev_8___repl2 (.Q (ENCR_DEV_prev_8___repl2), .D (
           nx15492z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_prev_8___repl3 (.Q (ENCR_DEV_prev_8___repl3), .D (
           nx15492z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_prev_8___repl4 (.Q (ENCR_DEV_prev_8___repl4), .D (
           nx15492z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_prev_8___repl5 (.Q (ENCR_DEV_prev_8___repl5), .D (
           nx15492z1), .CLK (CLK_int), .CLR (RST_int)) ;
    DFN1C0 ENCR_DEV_reg_prev_8___repl6 (.Q (ENCR_DEV_prev_8___repl6), .D (
           nx15492z1), .CLK (CLK_int), .CLR (RST_int)) ;
endmodule


module ram_dq_8_0 ( wr_data1, rd_data1, addr1, wr_clk1, rd_clk1, wr_ena1, 
                    rd_ena1, ena1, rst1, regce1, wr_data2, rd_data2, addr2, 
                    wr_clk2, rd_clk2, wr_ena2, rd_ena2, ena2, rst2, regce2, 
                    p_NOT_FIFO_DEV_rtlc5n43, p_RST_int, p_NOT_CONDITION_0_, 
                    p_WRITE, p_FIFO_DEV_rtlc_radd_N1_5___repl0, 
                    p_FIFO_DEV_rtlc_radd_N1_3___repl0, 
                    p_FIFO_DEV_rtlc_radd_N1_2___repl0, 
                    p_FIFO_DEV_rtlc_radd_N1_1___repl0, 
                    p_FIFO_DEV_rtlc_radd_N1_0___repl0 ) ;

    input [7:0]wr_data1 ;
    output [7:0]rd_data1 ;
    input [7:0]addr1 ;
    input wr_clk1 ;
    input rd_clk1 ;
    input wr_ena1 ;
    input rd_ena1 ;
    input ena1 ;
    input rst1 ;
    input regce1 ;
    input [7:0]wr_data2 ;
    output [7:0]rd_data2 ;
    input [7:0]addr2 ;
    input wr_clk2 ;
    input rd_clk2 ;
    input wr_ena2 ;
    input rd_ena2 ;
    input ena2 ;
    input rst2 ;
    input regce2 ;
    input p_NOT_FIFO_DEV_rtlc5n43 ;
    input p_RST_int ;
    input p_NOT_CONDITION_0_ ;
    input p_WRITE ;
    input p_FIFO_DEV_rtlc_radd_N1_5___repl0 ;
    input p_FIFO_DEV_rtlc_radd_N1_3___repl0 ;
    input p_FIFO_DEV_rtlc_radd_N1_2___repl0 ;
    input p_FIFO_DEV_rtlc_radd_N1_1___repl0 ;
    input p_FIFO_DEV_rtlc_radd_N1_0___repl0 ;

    wire nx9899z1, ena1_rename297, nx9899z2;
    wire [9:0] \$dummy ;




    RAM512X18 ix9899z43486 (.RD0 (rd_data2[0]), .RD1 (rd_data2[1]), .RD2 (
              rd_data2[2]), .RD3 (rd_data2[3]), .RD4 (rd_data2[4]), .RD5 (
              rd_data2[5]), .RD6 (rd_data2[6]), .RD7 (rd_data2[7]), .RD8 (
              \$dummy [0]), .RD9 (\$dummy [1]), .RD10 (\$dummy [2]), .RD11 (
              \$dummy [3]), .RD12 (\$dummy [4]), .RD13 (\$dummy [5]), .RD14 (
              \$dummy [6]), .RD15 (\$dummy [7]), .RD16 (\$dummy [8]), .RD17 (
              \$dummy [9]), .RADDR0 (p_FIFO_DEV_rtlc_radd_N1_0___repl0), .RADDR1 (
              p_FIFO_DEV_rtlc_radd_N1_1___repl0), .RADDR2 (
              p_FIFO_DEV_rtlc_radd_N1_2___repl0), .RADDR3 (
              p_FIFO_DEV_rtlc_radd_N1_3___repl0), .RADDR4 (addr2[4]), .RADDR5 (
              p_FIFO_DEV_rtlc_radd_N1_5___repl0), .RADDR6 (addr2[6]), .RADDR7 (
              addr2[7]), .RADDR8 (nx9899z1), .WADDR0 (addr1[0]), .WADDR1 (
              addr1[1]), .WADDR2 (addr1[2]), .WADDR3 (addr1[3]), .WADDR4 (
              addr1[4]), .WADDR5 (addr1[5]), .WADDR6 (addr1[6]), .WADDR7 (
              addr1[7]), .WADDR8 (nx9899z1), .WD0 (wr_data1[0]), .WD1 (
              wr_data1[1]), .WD2 (wr_data1[2]), .WD3 (wr_data1[3]), .WD4 (
              wr_data1[4]), .WD5 (wr_data1[5]), .WD6 (wr_data1[6]), .WD7 (
              wr_data1[7]), .WD8 (nx9899z1), .WD9 (nx9899z1), .WD10 (nx9899z1), 
              .WD11 (nx9899z1), .WD12 (nx9899z1), .WD13 (nx9899z1), .WD14 (
              nx9899z1), .WD15 (nx9899z1), .WD16 (nx9899z1), .WD17 (nx9899z1), .REN (
              nx9899z1), .WEN (nx9899z2), .RESET (ena1_rename297), .RW1 (
              nx9899z1), .RW0 (ena1_rename297), .WW1 (nx9899z1), .WW0 (
              ena1_rename297), .PIPE (nx9899z1), .RCLK (wr_clk1), .WCLK (wr_clk1
              )) ;
    GND ps_gnd (.Y (nx9899z1)) ;
    VCC ena1_rename301 (.Y (ena1_rename297)) ;
    NAND3 ix9899z24339 (.Y (nx9899z2), .A (p_RST_int), .B (p_NOT_CONDITION_0_), 
          .C (p_WRITE)) ;
endmodule


module mux_256_0 ( a, b, d, px994, px775, p_FIFO_DEV_rtlc_radd_N1_5___repl0, 
                   p_FIFO_DEV_rtlc_radd_N1_5___repl1, 
                   p_FIFO_DEV_rtlc_radd_N1_3___repl0, 
                   p_FIFO_DEV_rtlc_radd_N1_2___repl0, 
                   p_FIFO_DEV_rtlc_radd_N1_2___repl1, 
                   p_FIFO_DEV_rtlc_radd_N1_2___repl2, 
                   p_FIFO_DEV_rtlc_radd_N1_1___repl0, 
                   p_FIFO_DEV_rtlc_radd_N1_0___repl0 ) ;

    input [255:0]a ;
    input [255:0]b ;
    output d ;
    output px994 ;
    output px775 ;
    input p_FIFO_DEV_rtlc_radd_N1_5___repl0 ;
    input p_FIFO_DEV_rtlc_radd_N1_5___repl1 ;
    input p_FIFO_DEV_rtlc_radd_N1_3___repl0 ;
    input p_FIFO_DEV_rtlc_radd_N1_2___repl0 ;
    input p_FIFO_DEV_rtlc_radd_N1_2___repl1 ;
    input p_FIFO_DEV_rtlc_radd_N1_2___repl2 ;
    input p_FIFO_DEV_rtlc_radd_N1_1___repl0 ;
    input p_FIFO_DEV_rtlc_radd_N1_0___repl0 ;

    wire nx55823z65, nx14218z65, nx14218z97, nx14218z113, nx14218z121, 
         nx14218z125, nx14218z127, nx14218z114, nx14218z118, nx14218z120, 
         nx14218z98, nx14218z106, nx14218z110, nx14218z112, nx14218z99, 
         nx14218z103, nx14218z105, nx14218z66, nx14218z82, nx14218z90, 
         nx14218z94, nx14218z96, nx14218z83, nx14218z87, nx14218z89, nx14218z67, 
         nx14218z75, nx14218z79, nx14218z81, nx14218z68, nx14218z72, nx14218z74, 
         nx14218z122, nx14218z124, nx14218z115, nx14218z117, nx14218z107, 
         nx14218z109, nx14218z100, nx14218z102, nx14218z91, nx14218z93, 
         nx14218z84, nx14218z86, nx14218z76, nx14218z78, nx14218z69, nx14218z71, 
         nx14218z126, nx14218z119, nx14218z111, nx14218z104, nx14218z95, 
         nx14218z88, nx14218z80, nx14218z73, nx14218z123, nx14218z116, 
         nx14218z108, nx14218z101, nx14218z92, nx14218z85, nx14218z77, 
         nx14218z70, nx55823z97, nx55823z113, nx55823z121, nx55823z125, 
         nx55823z127, nx55823z114, nx55823z118, nx55823z120, nx55823z98, 
         nx55823z106, nx55823z110, nx55823z112, nx55823z99, nx55823z103, 
         nx55823z105, nx55823z66, nx55823z82, nx55823z90, nx55823z94, nx55823z96, 
         nx55823z83, nx55823z87, nx55823z89, nx55823z67, nx55823z75, nx55823z79, 
         nx55823z81, nx55823z68, nx55823z72, nx55823z74, nx55823z122, 
         nx55823z124, nx55823z115, nx55823z117, nx55823z107, nx55823z109, 
         nx55823z100, nx55823z102, nx55823z91, nx55823z93, nx55823z84, 
         nx55823z86, nx55823z76, nx55823z78, nx55823z69, nx55823z71, nx55823z126, 
         nx55823z119, nx55823z111, nx55823z104, nx55823z95, nx55823z88, 
         nx55823z80, nx55823z73, nx55823z123, nx55823z116, nx55823z108, 
         nx55823z101, nx55823z92, nx55823z85, nx55823z77, nx55823z70, nx55823z2, 
         nx55823z34, nx55823z50, nx55823z58, nx55823z62, nx55823z64, nx55823z59, 
         nx55823z61, nx55823z63, nx55823z60, nx55823z51, nx55823z55, nx55823z57, 
         nx55823z52, nx55823z54, nx55823z56, nx55823z53, nx55823z3, nx55823z19, 
         nx55823z27, nx55823z31, nx55823z33, nx55823z28, nx55823z30, nx55823z32, 
         nx55823z29, nx55823z20, nx55823z24, nx55823z26, nx55823z21, nx55823z23, 
         nx55823z25, nx55823z22, nx55823z35, nx55823z43, nx55823z47, nx55823z49, 
         nx55823z44, nx55823z46, nx55823z48, nx55823z45, nx55823z36, nx55823z40, 
         nx55823z42, nx55823z37, nx55823z39, nx55823z41, nx55823z38, nx55823z4, 
         nx55823z12, nx55823z16, nx55823z18, nx55823z13, nx55823z15, nx55823z17, 
         nx55823z14, nx55823z5, nx55823z9, nx55823z11, nx55823z6, nx55823z8, 
         nx55823z10, nx55823z7, nx14218z2, nx14218z34, nx14218z50, nx14218z58, 
         nx14218z62, nx14218z64, nx14218z59, nx14218z61, nx14218z51, nx14218z55, 
         nx14218z57, nx14218z52, nx14218z54, nx14218z35, nx14218z43, nx14218z47, 
         nx14218z49, nx14218z44, nx14218z46, nx14218z36, nx14218z40, nx14218z42, 
         nx14218z37, nx14218z39, nx14218z3, nx14218z19, nx14218z27, nx14218z31, 
         nx14218z33, nx14218z28, nx14218z30, nx14218z20, nx14218z24, nx14218z26, 
         nx14218z21, nx14218z23, nx14218z4, nx14218z12, nx14218z16, nx14218z18, 
         nx14218z13, nx14218z15, nx14218z5, nx14218z9, nx14218z11, nx14218z6, 
         nx14218z8, nx14218z63, nx14218z60, nx14218z56, nx14218z53, nx14218z48, 
         nx14218z45, nx14218z41, nx14218z38, nx14218z32, nx14218z29, nx14218z25, 
         nx14218z22, nx14218z17, nx14218z14, nx14218z10, nx14218z7;



    MX2 ix55823z14960 (.Y (nx55823z65), .A (nx55823z66), .S (b[3]), .B (
        nx55823z97)) ;
    MX2 ix14218z14960 (.Y (nx14218z65), .A (nx14218z66), .S (b[3]), .B (
        nx14218z97)) ;
    MX2 ix55823z14896 (.Y (px775), .A (nx55823z2), .S (b[6]), .B (nx55823z65)) ;
    MX2 ix14218z14992 (.Y (nx14218z97), .A (nx14218z98), .S (b[1]), .B (
        nx14218z113)) ;
    MX2 ix14218z15008 (.Y (nx14218z113), .A (nx14218z114), .S (b[0]), .B (
        nx14218z121)) ;
    MX2 ix14218z15016 (.Y (nx14218z121), .A (nx14218z122), .S (b[4]), .B (
        nx14218z125)) ;
    MX2 ix14218z15020 (.Y (nx14218z125), .A (nx14218z126), .S (b[5]), .B (
        nx14218z127)) ;
    MX2 ix14218z15022 (.Y (nx14218z127), .A (a[123]), .S (b[2]), .B (a[127])) ;
    MX2 ix14218z15009 (.Y (nx14218z114), .A (nx14218z115), .S (b[4]), .B (
        nx14218z118)) ;
    MX2 ix14218z15013 (.Y (nx14218z118), .A (nx14218z119), .S (b[5]), .B (
        nx14218z120)) ;
    MX2 ix14218z15015 (.Y (nx14218z120), .A (a[122]), .S (b[2]), .B (a[126])) ;
    MX2 ix14218z14993 (.Y (nx14218z98), .A (nx14218z99), .S (b[0]), .B (
        nx14218z106)) ;
    MX2 ix14218z15001 (.Y (nx14218z106), .A (nx14218z107), .S (b[4]), .B (
        nx14218z110)) ;
    MX2 ix14218z15005 (.Y (nx14218z110), .A (nx14218z111), .S (b[5]), .B (
        nx14218z112)) ;
    MX2 ix14218z15007 (.Y (nx14218z112), .A (a[121]), .S (b[2]), .B (a[125])) ;
    MX2 ix14218z14994 (.Y (nx14218z99), .A (nx14218z100), .S (b[4]), .B (
        nx14218z103)) ;
    MX2 ix14218z14998 (.Y (nx14218z103), .A (nx14218z104), .S (b[5]), .B (
        nx14218z105)) ;
    MX2 ix14218z15000 (.Y (nx14218z105), .A (a[120]), .S (b[2]), .B (a[124])) ;
    MX2 ix14218z14961 (.Y (nx14218z66), .A (nx14218z67), .S (b[1]), .B (
        nx14218z82)) ;
    MX2 ix14218z14977 (.Y (nx14218z82), .A (nx14218z83), .S (b[0]), .B (
        nx14218z90)) ;
    MX2 ix14218z14985 (.Y (nx14218z90), .A (nx14218z91), .S (b[4]), .B (
        nx14218z94)) ;
    MX2 ix14218z14989 (.Y (nx14218z94), .A (nx14218z95), .S (b[5]), .B (
        nx14218z96)) ;
    MX2 ix14218z14991 (.Y (nx14218z96), .A (a[115]), .S (b[2]), .B (a[119])) ;
    MX2 ix14218z14978 (.Y (nx14218z83), .A (nx14218z84), .S (b[4]), .B (
        nx14218z87)) ;
    MX2 ix14218z14982 (.Y (nx14218z87), .A (nx14218z88), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx14218z89)) ;
    MX2 ix14218z14984 (.Y (nx14218z89), .A (a[114]), .S (b[2]), .B (a[118])) ;
    MX2 ix14218z14962 (.Y (nx14218z67), .A (nx14218z68), .S (b[0]), .B (
        nx14218z75)) ;
    MX2 ix14218z14970 (.Y (nx14218z75), .A (nx14218z76), .S (b[4]), .B (
        nx14218z79)) ;
    MX2 ix14218z14974 (.Y (nx14218z79), .A (nx14218z80), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx14218z81)) ;
    MX2 ix14218z14976 (.Y (nx14218z81), .A (a[113]), .S (b[2]), .B (a[117])) ;
    MX2 ix14218z14963 (.Y (nx14218z68), .A (nx14218z69), .S (b[4]), .B (
        nx14218z72)) ;
    MX2 ix14218z14967 (.Y (nx14218z72), .A (nx14218z73), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx14218z74)) ;
    MX2 ix14218z14969 (.Y (nx14218z74), .A (a[112]), .S (b[2]), .B (a[116])) ;
    MX2 ix14218z15017 (.Y (nx14218z122), .A (nx14218z123), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx14218z124)) ;
    MX2 ix14218z15019 (.Y (nx14218z124), .A (a[107]), .S (b[2]), .B (a[111])) ;
    MX2 ix14218z15010 (.Y (nx14218z115), .A (nx14218z116), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx14218z117)) ;
    MX2 ix14218z15012 (.Y (nx14218z117), .A (a[106]), .S (b[2]), .B (a[110])) ;
    MX2 ix14218z15002 (.Y (nx14218z107), .A (nx14218z108), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx14218z109)) ;
    MX2 ix14218z15004 (.Y (nx14218z109), .A (a[105]), .S (b[2]), .B (a[109])) ;
    MX2 ix14218z14995 (.Y (nx14218z100), .A (nx14218z101), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx14218z102)) ;
    MX2 ix14218z14997 (.Y (nx14218z102), .A (a[104]), .S (b[2]), .B (a[108])) ;
    MX2 ix14218z14986 (.Y (nx14218z91), .A (nx14218z92), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx14218z93)) ;
    MX2 ix14218z14988 (.Y (nx14218z93), .A (a[99]), .S (b[2]), .B (a[103])) ;
    MX2 ix14218z14979 (.Y (nx14218z84), .A (nx14218z85), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx14218z86)) ;
    MX2 ix14218z14981 (.Y (nx14218z86), .A (a[98]), .S (b[2]), .B (a[102])) ;
    MX2 ix14218z14971 (.Y (nx14218z76), .A (nx14218z77), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx14218z78)) ;
    MX2 ix14218z14973 (.Y (nx14218z78), .A (a[97]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[101])) ;
    MX2 ix14218z14964 (.Y (nx14218z69), .A (nx14218z70), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx14218z71)) ;
    MX2 ix14218z14966 (.Y (nx14218z71), .A (a[96]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[100])) ;
    MX2 ix14218z15021 (.Y (nx14218z126), .A (a[91]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[95])) ;
    MX2 ix14218z15014 (.Y (nx14218z119), .A (a[90]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[94])) ;
    MX2 ix14218z15006 (.Y (nx14218z111), .A (a[89]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[93])) ;
    MX2 ix14218z14999 (.Y (nx14218z104), .A (a[88]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[92])) ;
    MX2 ix14218z14990 (.Y (nx14218z95), .A (a[83]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[87])) ;
    MX2 ix14218z14983 (.Y (nx14218z88), .A (a[82]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[86])) ;
    MX2 ix14218z14975 (.Y (nx14218z80), .A (a[81]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[85])) ;
    MX2 ix14218z14968 (.Y (nx14218z73), .A (a[80]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[84])) ;
    MX2 ix14218z15018 (.Y (nx14218z123), .A (a[75]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[79])) ;
    MX2 ix14218z15011 (.Y (nx14218z116), .A (a[74]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[78])) ;
    MX2 ix14218z15003 (.Y (nx14218z108), .A (a[73]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[77])) ;
    MX2 ix14218z14996 (.Y (nx14218z101), .A (a[72]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[76])) ;
    MX2 ix14218z14987 (.Y (nx14218z92), .A (a[67]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[71])) ;
    MX2 ix14218z14980 (.Y (nx14218z85), .A (a[66]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[70])) ;
    MX2 ix14218z14972 (.Y (nx14218z77), .A (a[65]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[69])) ;
    MX2 ix14218z14965 (.Y (nx14218z70), .A (a[64]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[68])) ;
    MX2 ix55823z14992 (.Y (nx55823z97), .A (nx55823z98), .S (b[1]), .B (
        nx55823z113)) ;
    MX2 ix55823z15008 (.Y (nx55823z113), .A (nx55823z114), .S (b[0]), .B (
        nx55823z121)) ;
    MX2 ix55823z15016 (.Y (nx55823z121), .A (nx55823z122), .S (b[4]), .B (
        nx55823z125)) ;
    MX2 ix55823z15020 (.Y (nx55823z125), .A (nx55823z126), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx55823z127)) ;
    MX2 ix55823z15022 (.Y (nx55823z127), .A (a[251]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[255])) ;
    MX2 ix55823z15009 (.Y (nx55823z114), .A (nx55823z115), .S (b[4]), .B (
        nx55823z118)) ;
    MX2 ix55823z15013 (.Y (nx55823z118), .A (nx55823z119), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx55823z120)) ;
    MX2 ix55823z15015 (.Y (nx55823z120), .A (a[250]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[254])) ;
    MX2 ix55823z14993 (.Y (nx55823z98), .A (nx55823z99), .S (
        p_FIFO_DEV_rtlc_radd_N1_0___repl0), .B (nx55823z106)) ;
    MX2 ix55823z15001 (.Y (nx55823z106), .A (nx55823z107), .S (b[4]), .B (
        nx55823z110)) ;
    MX2 ix55823z15005 (.Y (nx55823z110), .A (nx55823z111), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx55823z112)) ;
    MX2 ix55823z15007 (.Y (nx55823z112), .A (a[249]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[253])) ;
    MX2 ix55823z14994 (.Y (nx55823z99), .A (nx55823z100), .S (b[4]), .B (
        nx55823z103)) ;
    MX2 ix55823z14998 (.Y (nx55823z103), .A (nx55823z104), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx55823z105)) ;
    MX2 ix55823z15000 (.Y (nx55823z105), .A (a[248]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[252])) ;
    MX2 ix55823z14961 (.Y (nx55823z66), .A (nx55823z67), .S (b[1]), .B (
        nx55823z82)) ;
    MX2 ix55823z14977 (.Y (nx55823z82), .A (nx55823z83), .S (
        p_FIFO_DEV_rtlc_radd_N1_0___repl0), .B (nx55823z90)) ;
    MX2 ix55823z14985 (.Y (nx55823z90), .A (nx55823z91), .S (b[4]), .B (
        nx55823z94)) ;
    MX2 ix55823z14989 (.Y (nx55823z94), .A (nx55823z95), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx55823z96)) ;
    MX2 ix55823z14991 (.Y (nx55823z96), .A (a[243]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[247])) ;
    MX2 ix55823z14978 (.Y (nx55823z83), .A (nx55823z84), .S (b[4]), .B (
        nx55823z87)) ;
    MX2 ix55823z14982 (.Y (nx55823z87), .A (nx55823z88), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx55823z89)) ;
    MX2 ix55823z14984 (.Y (nx55823z89), .A (a[242]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl2), .B (a[246])) ;
    MX2 ix55823z14962 (.Y (nx55823z67), .A (nx55823z68), .S (
        p_FIFO_DEV_rtlc_radd_N1_0___repl0), .B (nx55823z75)) ;
    MX2 ix55823z14970 (.Y (nx55823z75), .A (nx55823z76), .S (b[4]), .B (
        nx55823z79)) ;
    MX2 ix55823z14974 (.Y (nx55823z79), .A (nx55823z80), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx55823z81)) ;
    MX2 ix55823z14976 (.Y (nx55823z81), .A (a[241]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[245])) ;
    MX2 ix55823z14963 (.Y (nx55823z68), .A (nx55823z69), .S (b[4]), .B (
        nx55823z72)) ;
    MX2 ix55823z14967 (.Y (nx55823z72), .A (nx55823z73), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx55823z74)) ;
    MX2 ix55823z14969 (.Y (nx55823z74), .A (a[240]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[244])) ;
    MX2 ix55823z15017 (.Y (nx55823z122), .A (nx55823z123), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx55823z124)) ;
    MX2 ix55823z15019 (.Y (nx55823z124), .A (a[235]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[239])) ;
    MX2 ix55823z15010 (.Y (nx55823z115), .A (nx55823z116), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx55823z117)) ;
    MX2 ix55823z15012 (.Y (nx55823z117), .A (a[234]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[238])) ;
    MX2 ix55823z15002 (.Y (nx55823z107), .A (nx55823z108), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx55823z109)) ;
    MX2 ix55823z15004 (.Y (nx55823z109), .A (a[233]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[237])) ;
    MX2 ix55823z14995 (.Y (nx55823z100), .A (nx55823z101), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx55823z102)) ;
    MX2 ix55823z14997 (.Y (nx55823z102), .A (a[232]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[236])) ;
    MX2 ix55823z14986 (.Y (nx55823z91), .A (nx55823z92), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl1), .B (nx55823z93)) ;
    MX2 ix55823z14988 (.Y (nx55823z93), .A (a[227]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[231])) ;
    MX2 ix55823z14979 (.Y (nx55823z84), .A (nx55823z85), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx55823z86)) ;
    MX2 ix55823z14981 (.Y (nx55823z86), .A (a[226]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[230])) ;
    MX2 ix55823z14971 (.Y (nx55823z76), .A (nx55823z77), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx55823z78)) ;
    MX2 ix55823z14973 (.Y (nx55823z78), .A (a[225]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[229])) ;
    MX2 ix55823z14964 (.Y (nx55823z69), .A (nx55823z70), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx55823z71)) ;
    MX2 ix55823z14966 (.Y (nx55823z71), .A (a[224]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[228])) ;
    MX2 ix55823z15021 (.Y (nx55823z126), .A (a[219]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[223])) ;
    MX2 ix55823z15014 (.Y (nx55823z119), .A (a[218]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[222])) ;
    MX2 ix55823z15006 (.Y (nx55823z111), .A (a[217]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[221])) ;
    MX2 ix55823z14999 (.Y (nx55823z104), .A (a[216]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[220])) ;
    MX2 ix55823z14990 (.Y (nx55823z95), .A (a[211]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[215])) ;
    MX2 ix55823z14983 (.Y (nx55823z88), .A (a[210]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[214])) ;
    MX2 ix55823z14975 (.Y (nx55823z80), .A (a[209]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[213])) ;
    MX2 ix55823z14968 (.Y (nx55823z73), .A (a[208]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[212])) ;
    MX2 ix55823z15018 (.Y (nx55823z123), .A (a[203]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[207])) ;
    MX2 ix55823z15011 (.Y (nx55823z116), .A (a[202]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[206])) ;
    MX2 ix55823z15003 (.Y (nx55823z108), .A (a[201]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[205])) ;
    MX2 ix55823z14996 (.Y (nx55823z101), .A (a[200]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[204])) ;
    MX2 ix55823z14987 (.Y (nx55823z92), .A (a[195]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[199])) ;
    MX2 ix55823z14980 (.Y (nx55823z85), .A (a[194]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl1), .B (a[198])) ;
    MX2 ix55823z14972 (.Y (nx55823z77), .A (a[193]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl0), .B (a[197])) ;
    MX2 ix55823z14965 (.Y (nx55823z70), .A (a[192]), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl0), .B (a[196])) ;
    MX2 ix55823z14897 (.Y (nx55823z2), .A (nx55823z3), .S (b[4]), .B (nx55823z34
        )) ;
    MX2 ix55823z14929 (.Y (nx55823z34), .A (nx55823z35), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx55823z50)) ;
    MX2 ix55823z14945 (.Y (nx55823z50), .A (nx55823z51), .S (b[3]), .B (
        nx55823z58)) ;
    MX2 ix55823z14953 (.Y (nx55823z58), .A (nx55823z59), .S (
        p_FIFO_DEV_rtlc_radd_N1_0___repl0), .B (nx55823z62)) ;
    MX2 ix55823z14957 (.Y (nx55823z62), .A (nx55823z63), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl0), .B (nx55823z64)) ;
    MX2 ix55823z14959 (.Y (nx55823z64), .A (a[189]), .S (b[1]), .B (a[191])) ;
    MX2 ix55823z14954 (.Y (nx55823z59), .A (nx55823z60), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl0), .B (nx55823z61)) ;
    MX2 ix55823z14956 (.Y (nx55823z61), .A (a[188]), .S (b[1]), .B (a[190])) ;
    MX2 ix55823z14958 (.Y (nx55823z63), .A (a[185]), .S (b[1]), .B (a[187])) ;
    MX2 ix55823z14955 (.Y (nx55823z60), .A (a[184]), .S (b[1]), .B (a[186])) ;
    MX2 ix55823z14946 (.Y (nx55823z51), .A (nx55823z52), .S (
        p_FIFO_DEV_rtlc_radd_N1_0___repl0), .B (nx55823z55)) ;
    MX2 ix55823z14950 (.Y (nx55823z55), .A (nx55823z56), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl0), .B (nx55823z57)) ;
    MX2 ix55823z14952 (.Y (nx55823z57), .A (a[181]), .S (b[1]), .B (a[183])) ;
    MX2 ix55823z14947 (.Y (nx55823z52), .A (nx55823z53), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl0), .B (nx55823z54)) ;
    MX2 ix55823z14949 (.Y (nx55823z54), .A (a[180]), .S (b[1]), .B (a[182])) ;
    MX2 ix55823z14951 (.Y (nx55823z56), .A (a[177]), .S (b[1]), .B (a[179])) ;
    MX2 ix55823z14948 (.Y (nx55823z53), .A (a[176]), .S (b[1]), .B (a[178])) ;
    MX2 ix55823z14898 (.Y (nx55823z3), .A (nx55823z4), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx55823z19)) ;
    MX2 ix55823z14914 (.Y (nx55823z19), .A (nx55823z20), .S (b[3]), .B (
        nx55823z27)) ;
    MX2 ix55823z14922 (.Y (nx55823z27), .A (nx55823z28), .S (
        p_FIFO_DEV_rtlc_radd_N1_0___repl0), .B (nx55823z31)) ;
    MX2 ix55823z14926 (.Y (nx55823z31), .A (nx55823z32), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl0), .B (nx55823z33)) ;
    MX2 ix55823z14928 (.Y (nx55823z33), .A (a[173]), .S (b[1]), .B (a[175])) ;
    MX2 ix55823z14923 (.Y (nx55823z28), .A (nx55823z29), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl0), .B (nx55823z30)) ;
    MX2 ix55823z14925 (.Y (nx55823z30), .A (a[172]), .S (b[1]), .B (a[174])) ;
    MX2 ix55823z14927 (.Y (nx55823z32), .A (a[169]), .S (b[1]), .B (a[171])) ;
    MX2 ix55823z14924 (.Y (nx55823z29), .A (a[168]), .S (b[1]), .B (a[170])) ;
    MX2 ix55823z14915 (.Y (nx55823z20), .A (nx55823z21), .S (
        p_FIFO_DEV_rtlc_radd_N1_0___repl0), .B (nx55823z24)) ;
    MX2 ix55823z14919 (.Y (nx55823z24), .A (nx55823z25), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl0), .B (nx55823z26)) ;
    MX2 ix55823z14921 (.Y (nx55823z26), .A (a[165]), .S (b[1]), .B (a[167])) ;
    MX2 ix55823z14916 (.Y (nx55823z21), .A (nx55823z22), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl0), .B (nx55823z23)) ;
    MX2 ix55823z14918 (.Y (nx55823z23), .A (a[164]), .S (b[1]), .B (a[166])) ;
    MX2 ix55823z14920 (.Y (nx55823z25), .A (a[161]), .S (b[1]), .B (a[163])) ;
    MX2 ix55823z14917 (.Y (nx55823z22), .A (a[160]), .S (b[1]), .B (a[162])) ;
    MX2 ix55823z14930 (.Y (nx55823z35), .A (nx55823z36), .S (b[3]), .B (
        nx55823z43)) ;
    MX2 ix55823z14938 (.Y (nx55823z43), .A (nx55823z44), .S (
        p_FIFO_DEV_rtlc_radd_N1_0___repl0), .B (nx55823z47)) ;
    MX2 ix55823z14942 (.Y (nx55823z47), .A (nx55823z48), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl0), .B (nx55823z49)) ;
    MX2 ix55823z14944 (.Y (nx55823z49), .A (a[157]), .S (
        p_FIFO_DEV_rtlc_radd_N1_1___repl0), .B (a[159])) ;
    MX2 ix55823z14939 (.Y (nx55823z44), .A (nx55823z45), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl0), .B (nx55823z46)) ;
    MX2 ix55823z14941 (.Y (nx55823z46), .A (a[156]), .S (
        p_FIFO_DEV_rtlc_radd_N1_1___repl0), .B (a[158])) ;
    MX2 ix55823z14943 (.Y (nx55823z48), .A (a[153]), .S (
        p_FIFO_DEV_rtlc_radd_N1_1___repl0), .B (a[155])) ;
    MX2 ix55823z14940 (.Y (nx55823z45), .A (a[152]), .S (
        p_FIFO_DEV_rtlc_radd_N1_1___repl0), .B (a[154])) ;
    MX2 ix55823z14931 (.Y (nx55823z36), .A (nx55823z37), .S (
        p_FIFO_DEV_rtlc_radd_N1_0___repl0), .B (nx55823z40)) ;
    MX2 ix55823z14935 (.Y (nx55823z40), .A (nx55823z41), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl0), .B (nx55823z42)) ;
    MX2 ix55823z14937 (.Y (nx55823z42), .A (a[149]), .S (
        p_FIFO_DEV_rtlc_radd_N1_1___repl0), .B (a[151])) ;
    MX2 ix55823z14932 (.Y (nx55823z37), .A (nx55823z38), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl0), .B (nx55823z39)) ;
    MX2 ix55823z14934 (.Y (nx55823z39), .A (a[148]), .S (
        p_FIFO_DEV_rtlc_radd_N1_1___repl0), .B (a[150])) ;
    MX2 ix55823z14936 (.Y (nx55823z41), .A (a[145]), .S (
        p_FIFO_DEV_rtlc_radd_N1_1___repl0), .B (a[147])) ;
    MX2 ix55823z14933 (.Y (nx55823z38), .A (a[144]), .S (
        p_FIFO_DEV_rtlc_radd_N1_1___repl0), .B (a[146])) ;
    MX2 ix55823z14899 (.Y (nx55823z4), .A (nx55823z5), .S (b[3]), .B (nx55823z12
        )) ;
    MX2 ix55823z14907 (.Y (nx55823z12), .A (nx55823z13), .S (
        p_FIFO_DEV_rtlc_radd_N1_0___repl0), .B (nx55823z16)) ;
    MX2 ix55823z14911 (.Y (nx55823z16), .A (nx55823z17), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl0), .B (nx55823z18)) ;
    MX2 ix55823z14913 (.Y (nx55823z18), .A (a[141]), .S (
        p_FIFO_DEV_rtlc_radd_N1_1___repl0), .B (a[143])) ;
    MX2 ix55823z14908 (.Y (nx55823z13), .A (nx55823z14), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl0), .B (nx55823z15)) ;
    MX2 ix55823z14910 (.Y (nx55823z15), .A (a[140]), .S (
        p_FIFO_DEV_rtlc_radd_N1_1___repl0), .B (a[142])) ;
    MX2 ix55823z14912 (.Y (nx55823z17), .A (a[137]), .S (
        p_FIFO_DEV_rtlc_radd_N1_1___repl0), .B (a[139])) ;
    MX2 ix55823z14909 (.Y (nx55823z14), .A (a[136]), .S (
        p_FIFO_DEV_rtlc_radd_N1_1___repl0), .B (a[138])) ;
    MX2 ix55823z14900 (.Y (nx55823z5), .A (nx55823z6), .S (
        p_FIFO_DEV_rtlc_radd_N1_0___repl0), .B (nx55823z9)) ;
    MX2 ix55823z14904 (.Y (nx55823z9), .A (nx55823z10), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl0), .B (nx55823z11)) ;
    MX2 ix55823z14906 (.Y (nx55823z11), .A (a[133]), .S (
        p_FIFO_DEV_rtlc_radd_N1_1___repl0), .B (a[135])) ;
    MX2 ix55823z14901 (.Y (nx55823z6), .A (nx55823z7), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl0), .B (nx55823z8)) ;
    MX2 ix55823z14903 (.Y (nx55823z8), .A (a[132]), .S (
        p_FIFO_DEV_rtlc_radd_N1_1___repl0), .B (a[134])) ;
    MX2 ix55823z14905 (.Y (nx55823z10), .A (a[129]), .S (
        p_FIFO_DEV_rtlc_radd_N1_1___repl0), .B (a[131])) ;
    MX2 ix55823z14902 (.Y (nx55823z7), .A (a[128]), .S (
        p_FIFO_DEV_rtlc_radd_N1_1___repl0), .B (a[130])) ;
    MX2 ix14218z14896 (.Y (px994), .A (nx14218z2), .S (b[6]), .B (nx14218z65)) ;
    MX2 ix14218z14897 (.Y (nx14218z2), .A (nx14218z3), .S (b[4]), .B (nx14218z34
        )) ;
    MX2 ix14218z14929 (.Y (nx14218z34), .A (nx14218z35), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl0), .B (nx14218z50)) ;
    MX2 ix14218z14945 (.Y (nx14218z50), .A (nx14218z51), .S (
        p_FIFO_DEV_rtlc_radd_N1_1___repl0), .B (nx14218z58)) ;
    MX2 ix14218z14953 (.Y (nx14218z58), .A (nx14218z59), .S (
        p_FIFO_DEV_rtlc_radd_N1_0___repl0), .B (nx14218z62)) ;
    MX2 ix14218z14957 (.Y (nx14218z62), .A (nx14218z63), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx14218z64)) ;
    MX2 ix14218z14959 (.Y (nx14218z64), .A (a[55]), .S (b[3]), .B (a[63])) ;
    MX2 ix14218z14954 (.Y (nx14218z59), .A (nx14218z60), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx14218z61)) ;
    MX2 ix14218z14956 (.Y (nx14218z61), .A (a[54]), .S (b[3]), .B (a[62])) ;
    MX2 ix14218z14946 (.Y (nx14218z51), .A (nx14218z52), .S (
        p_FIFO_DEV_rtlc_radd_N1_0___repl0), .B (nx14218z55)) ;
    MX2 ix14218z14950 (.Y (nx14218z55), .A (nx14218z56), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx14218z57)) ;
    MX2 ix14218z14952 (.Y (nx14218z57), .A (a[53]), .S (b[3]), .B (a[61])) ;
    MX2 ix14218z14947 (.Y (nx14218z52), .A (nx14218z53), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx14218z54)) ;
    MX2 ix14218z14949 (.Y (nx14218z54), .A (a[52]), .S (b[3]), .B (a[60])) ;
    MX2 ix14218z14930 (.Y (nx14218z35), .A (nx14218z36), .S (
        p_FIFO_DEV_rtlc_radd_N1_1___repl0), .B (nx14218z43)) ;
    MX2 ix14218z14938 (.Y (nx14218z43), .A (nx14218z44), .S (
        p_FIFO_DEV_rtlc_radd_N1_0___repl0), .B (nx14218z47)) ;
    MX2 ix14218z14942 (.Y (nx14218z47), .A (nx14218z48), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx14218z49)) ;
    MX2 ix14218z14944 (.Y (nx14218z49), .A (a[51]), .S (b[3]), .B (a[59])) ;
    MX2 ix14218z14939 (.Y (nx14218z44), .A (nx14218z45), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx14218z46)) ;
    MX2 ix14218z14941 (.Y (nx14218z46), .A (a[50]), .S (b[3]), .B (a[58])) ;
    MX2 ix14218z14931 (.Y (nx14218z36), .A (nx14218z37), .S (
        p_FIFO_DEV_rtlc_radd_N1_0___repl0), .B (nx14218z40)) ;
    MX2 ix14218z14935 (.Y (nx14218z40), .A (nx14218z41), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx14218z42)) ;
    MX2 ix14218z14937 (.Y (nx14218z42), .A (a[49]), .S (b[3]), .B (a[57])) ;
    MX2 ix14218z14932 (.Y (nx14218z37), .A (nx14218z38), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx14218z39)) ;
    MX2 ix14218z14934 (.Y (nx14218z39), .A (a[48]), .S (b[3]), .B (a[56])) ;
    MX2 ix14218z14898 (.Y (nx14218z3), .A (nx14218z4), .S (
        p_FIFO_DEV_rtlc_radd_N1_2___repl0), .B (nx14218z19)) ;
    MX2 ix14218z14914 (.Y (nx14218z19), .A (nx14218z20), .S (
        p_FIFO_DEV_rtlc_radd_N1_1___repl0), .B (nx14218z27)) ;
    MX2 ix14218z14922 (.Y (nx14218z27), .A (nx14218z28), .S (
        p_FIFO_DEV_rtlc_radd_N1_0___repl0), .B (nx14218z31)) ;
    MX2 ix14218z14926 (.Y (nx14218z31), .A (nx14218z32), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx14218z33)) ;
    MX2 ix14218z14928 (.Y (nx14218z33), .A (a[39]), .S (b[3]), .B (a[47])) ;
    MX2 ix14218z14923 (.Y (nx14218z28), .A (nx14218z29), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx14218z30)) ;
    MX2 ix14218z14925 (.Y (nx14218z30), .A (a[38]), .S (b[3]), .B (a[46])) ;
    MX2 ix14218z14915 (.Y (nx14218z20), .A (nx14218z21), .S (
        p_FIFO_DEV_rtlc_radd_N1_0___repl0), .B (nx14218z24)) ;
    MX2 ix14218z14919 (.Y (nx14218z24), .A (nx14218z25), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx14218z26)) ;
    MX2 ix14218z14921 (.Y (nx14218z26), .A (a[37]), .S (b[3]), .B (a[45])) ;
    MX2 ix14218z14916 (.Y (nx14218z21), .A (nx14218z22), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx14218z23)) ;
    MX2 ix14218z14918 (.Y (nx14218z23), .A (a[36]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[44])) ;
    MX2 ix14218z14899 (.Y (nx14218z4), .A (nx14218z5), .S (
        p_FIFO_DEV_rtlc_radd_N1_1___repl0), .B (nx14218z12)) ;
    MX2 ix14218z14907 (.Y (nx14218z12), .A (nx14218z13), .S (
        p_FIFO_DEV_rtlc_radd_N1_0___repl0), .B (nx14218z16)) ;
    MX2 ix14218z14911 (.Y (nx14218z16), .A (nx14218z17), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx14218z18)) ;
    MX2 ix14218z14913 (.Y (nx14218z18), .A (a[35]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[43])) ;
    MX2 ix14218z14908 (.Y (nx14218z13), .A (nx14218z14), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx14218z15)) ;
    MX2 ix14218z14910 (.Y (nx14218z15), .A (a[34]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[42])) ;
    MX2 ix14218z14900 (.Y (nx14218z5), .A (nx14218z6), .S (
        p_FIFO_DEV_rtlc_radd_N1_0___repl0), .B (nx14218z9)) ;
    MX2 ix14218z14904 (.Y (nx14218z9), .A (nx14218z10), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx14218z11)) ;
    MX2 ix14218z14906 (.Y (nx14218z11), .A (a[33]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[41])) ;
    MX2 ix14218z14901 (.Y (nx14218z6), .A (nx14218z7), .S (
        p_FIFO_DEV_rtlc_radd_N1_5___repl0), .B (nx14218z8)) ;
    MX2 ix14218z14903 (.Y (nx14218z8), .A (a[32]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[40])) ;
    MX2 ix14218z14958 (.Y (nx14218z63), .A (a[23]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[31])) ;
    MX2 ix14218z14955 (.Y (nx14218z60), .A (a[22]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[30])) ;
    MX2 ix14218z14951 (.Y (nx14218z56), .A (a[21]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[29])) ;
    MX2 ix14218z14948 (.Y (nx14218z53), .A (a[20]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[28])) ;
    MX2 ix14218z14943 (.Y (nx14218z48), .A (a[19]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[27])) ;
    MX2 ix14218z14940 (.Y (nx14218z45), .A (a[18]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[26])) ;
    MX2 ix14218z14936 (.Y (nx14218z41), .A (a[17]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[25])) ;
    MX2 ix14218z14933 (.Y (nx14218z38), .A (a[16]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[24])) ;
    MX2 ix14218z14927 (.Y (nx14218z32), .A (a[7]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[15])) ;
    MX2 ix14218z14924 (.Y (nx14218z29), .A (a[6]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[14])) ;
    MX2 ix14218z14920 (.Y (nx14218z25), .A (a[5]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[13])) ;
    MX2 ix14218z14917 (.Y (nx14218z22), .A (a[4]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[12])) ;
    MX2 ix14218z14912 (.Y (nx14218z17), .A (a[3]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[11])) ;
    MX2 ix14218z14909 (.Y (nx14218z14), .A (a[2]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[10])) ;
    MX2 ix14218z14905 (.Y (nx14218z10), .A (a[1]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[9])) ;
    MX2 ix14218z14902 (.Y (nx14218z7), .A (a[0]), .S (
        p_FIFO_DEV_rtlc_radd_N1_3___repl0), .B (a[8])) ;
endmodule


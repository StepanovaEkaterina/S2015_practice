`timescale 1 ns / 1 ns

program TLM_uart
();
endprogram
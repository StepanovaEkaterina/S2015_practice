module Trivium
(	input logic 			clk,
	input logic 			rst,
	input logic 			key,
	input logic 			[7:0] data,
	input logic 			strob_data,
	input logic 			strob_key,
	input logic 			[1:0] fifo_cnd,
	
	output logic 			[7:0] stream,
	output logic 			wt_sgn,
	output logic 			[7:0] sign_reg);

	logic [92:0] 			reg_str_1;
	logic [83:0] 			reg_str_2;
	logic [110:0] 			reg_str_3; 
	logic [79:0] 			vector=80'h00000000000000000000; //Вектор инициализации
	logic [0:7] 			t_1, t_2, t_3;
	logic [7:0]     		z;
			
	logic [11:0] 			cnt_init;//Счетчик инициализации
	logic [63:0] 			err_cnt; //2^64
	logic [6:0] 			key_cnt;  //Счетчик элементов ключа
	logic [8:0] 			encry_cnt; //Счетчик зашифрованных данных
			
	logic [7:0] 			data_reg; //Регистр входных данных
	logic [79:0] 			key_reg; //Регистр ключа шифрования
	logic					strob_data_tmp;
		
	enum logic [5:0] {NoKey, GetKey, KeyOK, Init, Moving_Secret, Secret_Ready, Error, Error_Key, Total_RST} nxt, prev;
/*Переприсвоение состояний*/
always_ff@(posedge clk, negedge rst)
begin
	if (!rst)
		prev<=NoKey;
	else
		prev<=nxt;
end
/*Безопасный приём данных*/
always_ff@(posedge clk, negedge rst)
begin
	if (!rst)
	begin
		strob_data_tmp<=0;
		data_reg<=0;
	end
	else
	begin
		strob_data_tmp<=strob_data;
		data_reg<=data;
	end
end
/*Определение состояния статусного регистра*/
always_ff@(posedge clk, negedge rst)
begin
	if (!rst)
		sign_reg<=8'b00000000;
	else
	begin
		unique case (prev)
		NoKey:
			sign_reg<=8'b00000000;
		GetKey:
			sign_reg<=8'b00000000;
		Moving_Secret:
			sign_reg<=8'b00000001;
		Secret_Ready:
			sign_reg<=8'b00000010;
		Error:
			sign_reg<=8'b00000100;
		Error_Key:
			sign_reg<=8'b00001000;
		Total_RST:
			sign_reg<=8'b00010000;
		default:
		    sign_reg<=8'b00000000;
		endcase
	end
end
/*Описание переходов конечного автомата*/
always_comb
begin
	unique case (prev)
	NoKey:
	begin
		if (strob_key)
			nxt=GetKey;
		else
			nxt=NoKey;
	end
	GetKey:
	begin
		/*if (strob_key)
			nxt=GetKey;
		else
			nxt=KeyOK;*/
		if (key_cnt<7'b1001111)
			if (strob_key)
				nxt=GetKey;
			else
				nxt=Error_Key;
		else if (strob_key)
				nxt=Error_Key;
			else
				nxt=KeyOK;
	end
	KeyOK:
	begin
		if (strob_key)
			nxt=GetKey;
		else
			nxt=Init;
	end
	Init:
	begin
		if (strob_key)
			nxt=Error_Key;
		else if (cnt_init<11'b10001111111)
				nxt=Init;
			else
				nxt=Moving_Secret;
	end
	Moving_Secret:
	begin
		if (strob_key)
			nxt=GetKey;
		else if (err_cnt>=2**64-1)
				nxt=Error;
			else if (encry_cnt == 8'b11111111)
					nxt=Secret_Ready;
				else
					nxt=Moving_Secret;
	end
	Secret_Ready:
	begin
		if (fifo_cnd==2'b00)
			nxt=Moving_Secret;
		else
			nxt=Secret_Ready;
	end
	Error:
	begin
		if (strob_data)
			nxt=Total_RST;
		else if (strob_key)
				nxt=GetKey;
			else
				nxt=Error;
	end
	Error_Key:
		nxt=NoKey;
	Total_RST:
		nxt=NoKey;
	default:
		nxt=NoKey;
	endcase
end
/*Получение ключа в разных состояниях автомата*/
always_ff@(posedge clk, negedge rst)
begin
	if(!rst)
	begin
		key_cnt<=0;
		key_reg<=0;
	end
	else
		unique case(prev)
		NoKey:
			key_reg<={key_reg[78:0],key};
		GetKey:
		begin
			if (key_cnt<7'b1010000)
			begin
				key_reg<={key_reg[78:0],key};
				key_cnt<=key_cnt+1;
			end
		else
			begin
				key_reg<=key_reg;
				key_cnt<=key_cnt;
			end
		end
		KeyOK:
		begin
			key_cnt<=0;
			if (strob_key)
				key_reg<={key_reg[78:0],key};
		end
		Moving_Secret:
		begin
			if (strob_key)
				key_reg<={key_reg[78:0],key};
		end
		Error:
		begin
			if (strob_key)
				key_reg<={key_reg[78:0],key};
		end
		Error_Key:
		begin
			key_cnt<=0;
			key_reg<=0;
		end
		Total_RST:
		begin
			key_cnt<=0;
			key_reg<=0;
		end
		default:
		begin
			key_cnt<=key_cnt;
			key_reg<=key_reg;
		end
		endcase
end
/*Блок шифрования и обновления счетчиков накопления и ошибок*/
always_ff@(posedge clk, negedge rst)
begin
  if (!rst)
  begin
	stream<=0;
	wt_sgn<=0;
	reg_str_1<=0;
	reg_str_2<=0;
	reg_str_3<=0;
	cnt_init<=0;
	err_cnt<=0;
	encry_cnt<=0;
  end
  else
  begin
	wt_sgn<=0;
	unique case(prev)
	GetKey:
	begin
		reg_str_1<=0;
		reg_str_2<=0;
		reg_str_3<=0;
	end
	KeyOK:
	begin
		reg_str_1[77:0]<=key_reg[79:2];
		reg_str_2[79:0]<=vector;
		reg_str_3[110:108]<=3'b111;
	end
	Init:
	begin
		reg_str_1<={reg_str_1[91:0], reg_str_3[65]^reg_str_3[110]^reg_str_3[108]&reg_str_3[109]^reg_str_1[68]};
		reg_str_2<={reg_str_2[82:0], reg_str_1[65]^reg_str_1[92] ^reg_str_1[90] &reg_str_1[91]^ reg_str_2[77]};
		reg_str_3<={reg_str_3[109:0],reg_str_2[68]^reg_str_2[83] ^reg_str_2[81] &reg_str_2[82]^ reg_str_3[86]};
		cnt_init<=cnt_init+1;
	end
	Moving_Secret:
	begin
	cnt_init<=0;
		if (strob_data_tmp)
		begin
			reg_str_1<={reg_str_1[84:0],t_3};
			reg_str_2<={reg_str_2[75:0],t_1};
			reg_str_3<={reg_str_3[102:0],t_2};
			stream<=data_reg^z;
			wt_sgn<=1;
			err_cnt<=err_cnt+1;
			encry_cnt<=encry_cnt+1;
		end
		else
		begin
			reg_str_1<=reg_str_1;
			reg_str_2<=reg_str_2;
			reg_str_3<=reg_str_3;
			wt_sgn<=0;
			stream<=0;
			err_cnt<=err_cnt;
			encry_cnt<=encry_cnt;
		end
	end
	Secret_Ready:
	begin
		encry_cnt<=0;
		stream<=0;
	end
	Total_RST:
	begin
		reg_str_1<=0;
		reg_str_2<=0;
		reg_str_3<=0;
		stream<=0;
		cnt_init<=0;
		err_cnt<=0;
		encry_cnt<=0;
	end
	default:
	begin
		stream<=stream;
		wt_sgn<=wt_sgn;
		reg_str_1<=reg_str_1;
		reg_str_2<=reg_str_2;
		reg_str_3<=reg_str_3;
		cnt_init<=cnt_init;
		err_cnt<=err_cnt;
		encry_cnt<=encry_cnt;
	end
  endcase
  end
end
/*Комбинационный блок для состояния шифрования*/
always_comb
begin
  for(int i=0;i<8;i++)
    begin
      z[i]=reg_str_1[65-i]^reg_str_1[92-i]^reg_str_2[68-i]^reg_str_2[83-i]^reg_str_3[65-i]^reg_str_3[110-i];
      t_1[i]=reg_str_1[65-i]^reg_str_1[92-i]^ reg_str_1[90-i]& reg_str_1[91-i]^ reg_str_2[77-i];
      t_2[i]=reg_str_2[68-i]^reg_str_2[83-i]^ reg_str_2[81-i]& reg_str_2[82-i]^ reg_str_3[86-i];
      t_3[i]=reg_str_3[65-i]^reg_str_3[110-i]^reg_str_3[108-i]&reg_str_3[109-i]^reg_str_1[68-i];
    end
end
endmodule